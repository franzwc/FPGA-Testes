//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2014 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_0_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_0_upstream_module (
                                                                                           // inputs:
                                                                                            clear_fifo,
                                                                                            clk,
                                                                                            data_in,
                                                                                            read,
                                                                                            reset_n,
                                                                                            sync_reset,
                                                                                            write,

                                                                                           // outputs:
                                                                                            data_out,
                                                                                            empty,
                                                                                            fifo_contains_ones_n,
                                                                                            full
                                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_0_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_0_upstream_readdata,
                                                   Medipix_sopc_burst_0_upstream_readdatavalid,
                                                   Medipix_sopc_burst_0_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_instruction_master_address_to_slave,
                                                   cpu_linux_instruction_master_burstcount,
                                                   cpu_linux_instruction_master_latency_counter,
                                                   cpu_linux_instruction_master_read,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_0_upstream_address,
                                                   Medipix_sopc_burst_0_upstream_byteaddress,
                                                   Medipix_sopc_burst_0_upstream_byteenable,
                                                   Medipix_sopc_burst_0_upstream_debugaccess,
                                                   Medipix_sopc_burst_0_upstream_read,
                                                   Medipix_sopc_burst_0_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_0_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_0_upstream_write,
                                                   cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream,
                                                   cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register,
                                                   cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream,
                                                   d1_Medipix_sopc_burst_0_upstream_end_xfer
                                                )
;

  output  [ 10: 0] Medipix_sopc_burst_0_upstream_address;
  output  [ 12: 0] Medipix_sopc_burst_0_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_0_upstream_byteenable;
  output           Medipix_sopc_burst_0_upstream_debugaccess;
  output           Medipix_sopc_burst_0_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_0_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_0_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_0_upstream_write;
  output           cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream;
  output           cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream;
  output           cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream;
  output           cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register;
  output           cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream;
  output           d1_Medipix_sopc_burst_0_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_0_upstream_readdata;
  input            Medipix_sopc_burst_0_upstream_readdatavalid;
  input            Medipix_sopc_burst_0_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_instruction_master_address_to_slave;
  input   [  3: 0] cpu_linux_instruction_master_burstcount;
  input            cpu_linux_instruction_master_latency_counter;
  input            cpu_linux_instruction_master_read;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register;
  input            reset_n;

  wire    [ 10: 0] Medipix_sopc_burst_0_upstream_address;
  wire             Medipix_sopc_burst_0_upstream_allgrants;
  wire             Medipix_sopc_burst_0_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_0_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_0_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_0_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_0_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_arb_share_set_values;
  wire             Medipix_sopc_burst_0_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_0_upstream_begins_xfer;
  wire             Medipix_sopc_burst_0_upstream_burstcount_fifo_empty;
  wire    [ 12: 0] Medipix_sopc_burst_0_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_0_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_0_upstream_debugaccess;
  wire             Medipix_sopc_burst_0_upstream_end_xfer;
  wire             Medipix_sopc_burst_0_upstream_firsttransfer;
  wire             Medipix_sopc_burst_0_upstream_grant_vector;
  wire             Medipix_sopc_burst_0_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_0_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_0_upstream_load_fifo;
  wire             Medipix_sopc_burst_0_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_0_upstream_move_on_to_next_transaction;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_next_burst_count;
  wire             Medipix_sopc_burst_0_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_0_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_0_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_0_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_0_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_0_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_0_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_0_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_0_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_0_upstream_waits_for_read;
  wire             Medipix_sopc_burst_0_upstream_waits_for_write;
  wire             Medipix_sopc_burst_0_upstream_write;
  wire             cpu_linux_instruction_master_arbiterlock;
  wire             cpu_linux_instruction_master_arbiterlock2;
  wire             cpu_linux_instruction_master_continuerequest;
  wire             cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_rdv_fifo_output_from_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register;
  wire             cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_0_upstream;
  reg              d1_Medipix_sopc_burst_0_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_0_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_0_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_0_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_0_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream));
  //assign Medipix_sopc_burst_0_upstream_readdata_from_sa = Medipix_sopc_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_readdata_from_sa = Medipix_sopc_burst_0_upstream_readdata;

  assign cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream = (({cpu_linux_instruction_master_address_to_slave[27 : 11] , 11'b0} == 28'h8003800) & (cpu_linux_instruction_master_read)) & cpu_linux_instruction_master_read;
  //assign Medipix_sopc_burst_0_upstream_waitrequest_from_sa = Medipix_sopc_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_waitrequest_from_sa = Medipix_sopc_burst_0_upstream_waitrequest;

  //assign Medipix_sopc_burst_0_upstream_readdatavalid_from_sa = Medipix_sopc_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_readdatavalid_from_sa = Medipix_sopc_burst_0_upstream_readdatavalid;

  //Medipix_sopc_burst_0_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_arb_share_set_values = 1;

  //Medipix_sopc_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_any_bursting_master_saved_grant = cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_0_upstream;

  //Medipix_sopc_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_arb_share_counter_next_value = Medipix_sopc_burst_0_upstream_firsttransfer ? (Medipix_sopc_burst_0_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_0_upstream_arb_share_counter ? (Medipix_sopc_burst_0_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_0_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_allgrants = |Medipix_sopc_burst_0_upstream_grant_vector;

  //Medipix_sopc_burst_0_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_end_xfer = ~(Medipix_sopc_burst_0_upstream_waits_for_read | Medipix_sopc_burst_0_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream = Medipix_sopc_burst_0_upstream_end_xfer & (~Medipix_sopc_burst_0_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream & Medipix_sopc_burst_0_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream & ~Medipix_sopc_burst_0_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_0_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_0_upstream_arb_counter_enable)
          Medipix_sopc_burst_0_upstream_arb_share_counter <= Medipix_sopc_burst_0_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_0_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_0_upstream & ~Medipix_sopc_burst_0_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_0_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_0_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/instruction_master Medipix_sopc_burst_0/upstream arbiterlock, which is an e_assign
  assign cpu_linux_instruction_master_arbiterlock = Medipix_sopc_burst_0_upstream_slavearbiterlockenable & cpu_linux_instruction_master_continuerequest;

  //Medipix_sopc_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_0_upstream_arb_share_counter_next_value;

  //cpu_linux/instruction_master Medipix_sopc_burst_0/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_instruction_master_arbiterlock2 = Medipix_sopc_burst_0_upstream_slavearbiterlockenable2 & cpu_linux_instruction_master_continuerequest;

  //Medipix_sopc_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_any_continuerequest = 1;

  //cpu_linux_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_instruction_master_continuerequest = 1;

  assign cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream = cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream & ~((cpu_linux_instruction_master_read & ((cpu_linux_instruction_master_latency_counter != 0) | (1 < cpu_linux_instruction_master_latency_counter) | (|cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register) | (|cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_move_on_to_next_transaction = Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_0_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_0_upstream, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_selected_burstcount = (cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream)? cpu_linux_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_0_upstream_module burstcount_fifo_for_Medipix_sopc_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_0_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_0_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_0_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read & Medipix_sopc_burst_0_upstream_load_fifo & ~(Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_0_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_0_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_current_burst_minus_one = Medipix_sopc_burst_0_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_0_upstream, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read) & ~Medipix_sopc_burst_0_upstream_load_fifo))? Medipix_sopc_burst_0_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read & Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_0_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_0_upstream_selected_burstcount :
    (Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_0_upstream_transaction_burst_count :
    Medipix_sopc_burst_0_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_0_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_0_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_0_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read)))
          Medipix_sopc_burst_0_upstream_current_burst <= Medipix_sopc_burst_0_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_0_upstream_load_fifo = (~Medipix_sopc_burst_0_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read) & Medipix_sopc_burst_0_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_0_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read) & ~Medipix_sopc_burst_0_upstream_load_fifo | Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_0_upstream_load_fifo <= p0_Medipix_sopc_burst_0_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_0_upstream, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_0_upstream_current_burst_minus_one) & Medipix_sopc_burst_0_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_0_upstream_module rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream),
      .data_out             (cpu_linux_instruction_master_rdv_fifo_output_from_Medipix_sopc_burst_0_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_0_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_0_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_0_upstream_waits_for_read)
    );

  assign cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register = ~cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_0_upstream;
  //local readdatavalid cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream, which is an e_mux
  assign cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream = Medipix_sopc_burst_0_upstream_readdatavalid_from_sa;

  //byteaddress mux for Medipix_sopc_burst_0/upstream, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_byteaddress = cpu_linux_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream = cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream;

  //cpu_linux/instruction_master saved-grant Medipix_sopc_burst_0/upstream, which is an e_assign
  assign cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_0_upstream = cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream;

  //allow new arb cycle for Medipix_sopc_burst_0/upstream, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_0_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_0_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_firsttransfer = Medipix_sopc_burst_0_upstream_begins_xfer ? Medipix_sopc_burst_0_upstream_unreg_firsttransfer : Medipix_sopc_burst_0_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_0_upstream_slavearbiterlockenable & Medipix_sopc_burst_0_upstream_any_continuerequest);

  //Medipix_sopc_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_0_upstream_begins_xfer)
          Medipix_sopc_burst_0_upstream_reg_firsttransfer <= Medipix_sopc_burst_0_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_beginbursttransfer_internal = Medipix_sopc_burst_0_upstream_begins_xfer;

  //Medipix_sopc_burst_0_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_read = cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream & cpu_linux_instruction_master_read;

  //Medipix_sopc_burst_0_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_write = 0;

  //Medipix_sopc_burst_0_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_address = cpu_linux_instruction_master_address_to_slave;

  //d1_Medipix_sopc_burst_0_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_0_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_0_upstream_end_xfer <= Medipix_sopc_burst_0_upstream_end_xfer;
    end


  //Medipix_sopc_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_waits_for_read = Medipix_sopc_burst_0_upstream_in_a_read_cycle & Medipix_sopc_burst_0_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_in_a_read_cycle = cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream & cpu_linux_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_0_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_waits_for_write = Medipix_sopc_burst_0_upstream_in_a_write_cycle & Medipix_sopc_burst_0_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_0_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_0_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_0_upstream_counter = 0;
  //Medipix_sopc_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_0_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_0/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream && (cpu_linux_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/instruction_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_0/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_0_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_0_downstream_address,
                                                     Medipix_sopc_burst_0_downstream_burstcount,
                                                     Medipix_sopc_burst_0_downstream_byteenable,
                                                     Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_0_downstream_read,
                                                     Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_0_downstream_write,
                                                     Medipix_sopc_burst_0_downstream_writedata,
                                                     clk,
                                                     cpu_linux_jtag_debug_module_readdata_from_sa,
                                                     d1_cpu_linux_jtag_debug_module_end_xfer,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_0_downstream_address_to_slave,
                                                     Medipix_sopc_burst_0_downstream_latency_counter,
                                                     Medipix_sopc_burst_0_downstream_readdata,
                                                     Medipix_sopc_burst_0_downstream_readdatavalid,
                                                     Medipix_sopc_burst_0_downstream_reset_n,
                                                     Medipix_sopc_burst_0_downstream_waitrequest
                                                  )
;

  output  [ 10: 0] Medipix_sopc_burst_0_downstream_address_to_slave;
  output           Medipix_sopc_burst_0_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_0_downstream_readdata;
  output           Medipix_sopc_burst_0_downstream_readdatavalid;
  output           Medipix_sopc_burst_0_downstream_reset_n;
  output           Medipix_sopc_burst_0_downstream_waitrequest;
  input   [ 10: 0] Medipix_sopc_burst_0_downstream_address;
  input            Medipix_sopc_burst_0_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_0_downstream_byteenable;
  input            Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_0_downstream_read;
  input            Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_0_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_0_downstream_writedata;
  input            clk;
  input   [ 31: 0] cpu_linux_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_linux_jtag_debug_module_end_xfer;
  input            reset_n;

  reg     [ 10: 0] Medipix_sopc_burst_0_downstream_address_last_time;
  wire    [ 10: 0] Medipix_sopc_burst_0_downstream_address_to_slave;
  reg              Medipix_sopc_burst_0_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_0_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_0_downstream_is_granted_some_slave;
  reg              Medipix_sopc_burst_0_downstream_latency_counter;
  reg              Medipix_sopc_burst_0_downstream_read_but_no_slave_selected;
  reg              Medipix_sopc_burst_0_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_0_downstream_readdata;
  wire             Medipix_sopc_burst_0_downstream_readdatavalid;
  wire             Medipix_sopc_burst_0_downstream_reset_n;
  wire             Medipix_sopc_burst_0_downstream_run;
  wire             Medipix_sopc_burst_0_downstream_waitrequest;
  reg              Medipix_sopc_burst_0_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_0_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_Medipix_sopc_burst_0_downstream_latency_counter;
  wire             pre_flush_Medipix_sopc_burst_0_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module) & (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module) & ((~Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_0_downstream_read | (1 & ~d1_cpu_linux_jtag_debug_module_end_xfer & Medipix_sopc_burst_0_downstream_read))) & ((~Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_0_downstream_write | (1 & Medipix_sopc_burst_0_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_0_downstream_address_to_slave = Medipix_sopc_burst_0_downstream_address;

  //Medipix_sopc_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_read_but_no_slave_selected <= 0;
      else 
        Medipix_sopc_burst_0_downstream_read_but_no_slave_selected <= Medipix_sopc_burst_0_downstream_read & Medipix_sopc_burst_0_downstream_run & ~Medipix_sopc_burst_0_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign Medipix_sopc_burst_0_downstream_is_granted_some_slave = Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_0_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_0_downstream_readdatavalid = Medipix_sopc_burst_0_downstream_read_but_no_slave_selected |
    pre_flush_Medipix_sopc_burst_0_downstream_readdatavalid |
    Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module;

  //Medipix_sopc_burst_0/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_0_downstream_readdata = cpu_linux_jtag_debug_module_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_waitrequest = ~Medipix_sopc_burst_0_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_latency_counter <= 0;
      else 
        Medipix_sopc_burst_0_downstream_latency_counter <= p1_Medipix_sopc_burst_0_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_Medipix_sopc_burst_0_downstream_latency_counter = ((Medipix_sopc_burst_0_downstream_run & Medipix_sopc_burst_0_downstream_read))? latency_load_value :
    (Medipix_sopc_burst_0_downstream_latency_counter)? Medipix_sopc_burst_0_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //Medipix_sopc_burst_0_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_0_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_0_downstream_address_last_time <= Medipix_sopc_burst_0_downstream_address;
    end


  //Medipix_sopc_burst_0/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_0_downstream_waitrequest & (Medipix_sopc_burst_0_downstream_read | Medipix_sopc_burst_0_downstream_write);
    end


  //Medipix_sopc_burst_0_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_0_downstream_address != Medipix_sopc_burst_0_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_0_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_0_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_0_downstream_burstcount_last_time <= Medipix_sopc_burst_0_downstream_burstcount;
    end


  //Medipix_sopc_burst_0_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_0_downstream_burstcount != Medipix_sopc_burst_0_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_0_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_0_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_0_downstream_byteenable_last_time <= Medipix_sopc_burst_0_downstream_byteenable;
    end


  //Medipix_sopc_burst_0_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_0_downstream_byteenable != Medipix_sopc_burst_0_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_0_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_0_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_0_downstream_read_last_time <= Medipix_sopc_burst_0_downstream_read;
    end


  //Medipix_sopc_burst_0_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_0_downstream_read != Medipix_sopc_burst_0_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_0_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_0_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_0_downstream_write_last_time <= Medipix_sopc_burst_0_downstream_write;
    end


  //Medipix_sopc_burst_0_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_0_downstream_write != Medipix_sopc_burst_0_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_0_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_0_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_0_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_0_downstream_writedata_last_time <= Medipix_sopc_burst_0_downstream_writedata;
    end


  //Medipix_sopc_burst_0_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_0_downstream_writedata != Medipix_sopc_burst_0_downstream_writedata_last_time) & Medipix_sopc_burst_0_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_0_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_1_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_1_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_1_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_1_upstream_readdata,
                                                   Medipix_sopc_burst_1_upstream_readdatavalid,
                                                   Medipix_sopc_burst_1_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_1_upstream_address,
                                                   Medipix_sopc_burst_1_upstream_burstcount,
                                                   Medipix_sopc_burst_1_upstream_byteaddress,
                                                   Medipix_sopc_burst_1_upstream_byteenable,
                                                   Medipix_sopc_burst_1_upstream_debugaccess,
                                                   Medipix_sopc_burst_1_upstream_read,
                                                   Medipix_sopc_burst_1_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_1_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_1_upstream_write,
                                                   Medipix_sopc_burst_1_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream,
                                                   d1_Medipix_sopc_burst_1_upstream_end_xfer
                                                )
;

  output  [ 10: 0] Medipix_sopc_burst_1_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_1_upstream_burstcount;
  output  [ 12: 0] Medipix_sopc_burst_1_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_1_upstream_byteenable;
  output           Medipix_sopc_burst_1_upstream_debugaccess;
  output           Medipix_sopc_burst_1_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_1_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_1_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_1_upstream_write;
  output  [ 31: 0] Medipix_sopc_burst_1_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream;
  output           d1_Medipix_sopc_burst_1_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_1_upstream_readdata;
  input            Medipix_sopc_burst_1_upstream_readdatavalid;
  input            Medipix_sopc_burst_1_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [ 10: 0] Medipix_sopc_burst_1_upstream_address;
  wire             Medipix_sopc_burst_1_upstream_allgrants;
  wire             Medipix_sopc_burst_1_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_1_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_1_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_1_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_1_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_1_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_1_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_1_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_burstcount;
  wire             Medipix_sopc_burst_1_upstream_burstcount_fifo_empty;
  wire    [ 12: 0] Medipix_sopc_burst_1_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_1_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_1_upstream_debugaccess;
  wire             Medipix_sopc_burst_1_upstream_end_xfer;
  wire             Medipix_sopc_burst_1_upstream_firsttransfer;
  wire             Medipix_sopc_burst_1_upstream_grant_vector;
  wire             Medipix_sopc_burst_1_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_1_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_1_upstream_load_fifo;
  wire             Medipix_sopc_burst_1_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_1_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_1_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_next_burst_count;
  wire             Medipix_sopc_burst_1_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_1_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_1_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_1_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_1_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_1_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_1_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_1_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_1_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_1_upstream_waits_for_read;
  wire             Medipix_sopc_burst_1_upstream_waits_for_write;
  wire             Medipix_sopc_burst_1_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_1_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_1_upstream;
  reg              d1_Medipix_sopc_burst_1_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_1_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_1_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_1_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_1_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream));
  //assign Medipix_sopc_burst_1_upstream_readdata_from_sa = Medipix_sopc_burst_1_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_readdata_from_sa = Medipix_sopc_burst_1_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream = ({cpu_linux_data_master_address_to_slave[27 : 11] , 11'b0} == 28'h8003800) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_1_upstream_waitrequest_from_sa = Medipix_sopc_burst_1_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_waitrequest_from_sa = Medipix_sopc_burst_1_upstream_waitrequest;

  //assign Medipix_sopc_burst_1_upstream_readdatavalid_from_sa = Medipix_sopc_burst_1_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_readdatavalid_from_sa = Medipix_sopc_burst_1_upstream_readdatavalid;

  //Medipix_sopc_burst_1_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_1_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_1_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_1_upstream;

  //Medipix_sopc_burst_1_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_arb_share_counter_next_value = Medipix_sopc_burst_1_upstream_firsttransfer ? (Medipix_sopc_burst_1_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_1_upstream_arb_share_counter ? (Medipix_sopc_burst_1_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_1_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_allgrants = |Medipix_sopc_burst_1_upstream_grant_vector;

  //Medipix_sopc_burst_1_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_end_xfer = ~(Medipix_sopc_burst_1_upstream_waits_for_read | Medipix_sopc_burst_1_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream = Medipix_sopc_burst_1_upstream_end_xfer & (~Medipix_sopc_burst_1_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_1_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream & Medipix_sopc_burst_1_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream & ~Medipix_sopc_burst_1_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_1_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_1_upstream_arb_counter_enable)
          Medipix_sopc_burst_1_upstream_arb_share_counter <= Medipix_sopc_burst_1_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_1_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_1_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_1_upstream & ~Medipix_sopc_burst_1_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_1_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_1_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_1/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_1_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_1_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_1_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_1/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_1_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_1_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_1_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_move_on_to_next_transaction = Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_1_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_1_upstream, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_1_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_1_upstream_module burstcount_fifo_for_Medipix_sopc_burst_1_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_1_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_1_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_1_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read & Medipix_sopc_burst_1_upstream_load_fifo & ~(Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_1_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_1_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_current_burst_minus_one = Medipix_sopc_burst_1_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_1_upstream, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read) & ~Medipix_sopc_burst_1_upstream_load_fifo))? Medipix_sopc_burst_1_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read & Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_1_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_1_upstream_selected_burstcount :
    (Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_1_upstream_transaction_burst_count :
    Medipix_sopc_burst_1_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_1_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_1_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_1_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read)))
          Medipix_sopc_burst_1_upstream_current_burst <= Medipix_sopc_burst_1_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_1_upstream_load_fifo = (~Medipix_sopc_burst_1_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read) & Medipix_sopc_burst_1_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_1_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read) & ~Medipix_sopc_burst_1_upstream_load_fifo | Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_1_upstream_load_fifo <= p0_Medipix_sopc_burst_1_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_1_upstream, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_1_upstream_current_burst_minus_one) & Medipix_sopc_burst_1_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_1_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_1_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_1_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_1_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_1_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_1_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_1_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_1_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream = Medipix_sopc_burst_1_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_1_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_1/upstream, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_1/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_1_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream;

  //allow new arb cycle for Medipix_sopc_burst_1/upstream, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_1_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_1_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_1_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_firsttransfer = Medipix_sopc_burst_1_upstream_begins_xfer ? Medipix_sopc_burst_1_upstream_unreg_firsttransfer : Medipix_sopc_burst_1_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_1_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_1_upstream_slavearbiterlockenable & Medipix_sopc_burst_1_upstream_any_continuerequest);

  //Medipix_sopc_burst_1_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_1_upstream_begins_xfer)
          Medipix_sopc_burst_1_upstream_reg_firsttransfer <= Medipix_sopc_burst_1_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_1_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_1_upstream_write) && (Medipix_sopc_burst_1_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_1_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_1_upstream_read) && (Medipix_sopc_burst_1_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_1_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_1_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_1_upstream_begins_xfer)
          Medipix_sopc_burst_1_upstream_bbt_burstcounter <= Medipix_sopc_burst_1_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_1_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_beginbursttransfer_internal = Medipix_sopc_burst_1_upstream_begins_xfer & (Medipix_sopc_burst_1_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_1_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_1_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream & cpu_linux_data_master_write;

  //Medipix_sopc_burst_1_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_address = cpu_linux_data_master_address_to_slave;

  //d1_Medipix_sopc_burst_1_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_1_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_1_upstream_end_xfer <= Medipix_sopc_burst_1_upstream_end_xfer;
    end


  //Medipix_sopc_burst_1_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_waits_for_read = Medipix_sopc_burst_1_upstream_in_a_read_cycle & Medipix_sopc_burst_1_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_1_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_1_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_1_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_waits_for_write = Medipix_sopc_burst_1_upstream_in_a_write_cycle & Medipix_sopc_burst_1_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_1_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_1_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_1_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_1_upstream_counter = 0;
  //Medipix_sopc_burst_1_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_1_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_1/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_1/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_1_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_1_downstream_address,
                                                     Medipix_sopc_burst_1_downstream_burstcount,
                                                     Medipix_sopc_burst_1_downstream_byteenable,
                                                     Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_1_downstream_read,
                                                     Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module,
                                                     Medipix_sopc_burst_1_downstream_write,
                                                     Medipix_sopc_burst_1_downstream_writedata,
                                                     clk,
                                                     cpu_linux_jtag_debug_module_readdata_from_sa,
                                                     d1_cpu_linux_jtag_debug_module_end_xfer,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_1_downstream_address_to_slave,
                                                     Medipix_sopc_burst_1_downstream_latency_counter,
                                                     Medipix_sopc_burst_1_downstream_readdata,
                                                     Medipix_sopc_burst_1_downstream_readdatavalid,
                                                     Medipix_sopc_burst_1_downstream_reset_n,
                                                     Medipix_sopc_burst_1_downstream_waitrequest
                                                  )
;

  output  [ 10: 0] Medipix_sopc_burst_1_downstream_address_to_slave;
  output           Medipix_sopc_burst_1_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_1_downstream_readdata;
  output           Medipix_sopc_burst_1_downstream_readdatavalid;
  output           Medipix_sopc_burst_1_downstream_reset_n;
  output           Medipix_sopc_burst_1_downstream_waitrequest;
  input   [ 10: 0] Medipix_sopc_burst_1_downstream_address;
  input            Medipix_sopc_burst_1_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_1_downstream_byteenable;
  input            Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_1_downstream_read;
  input            Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module;
  input            Medipix_sopc_burst_1_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_1_downstream_writedata;
  input            clk;
  input   [ 31: 0] cpu_linux_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_linux_jtag_debug_module_end_xfer;
  input            reset_n;

  reg     [ 10: 0] Medipix_sopc_burst_1_downstream_address_last_time;
  wire    [ 10: 0] Medipix_sopc_burst_1_downstream_address_to_slave;
  reg              Medipix_sopc_burst_1_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_1_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_1_downstream_is_granted_some_slave;
  reg              Medipix_sopc_burst_1_downstream_latency_counter;
  reg              Medipix_sopc_burst_1_downstream_read_but_no_slave_selected;
  reg              Medipix_sopc_burst_1_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_1_downstream_readdata;
  wire             Medipix_sopc_burst_1_downstream_readdatavalid;
  wire             Medipix_sopc_burst_1_downstream_reset_n;
  wire             Medipix_sopc_burst_1_downstream_run;
  wire             Medipix_sopc_burst_1_downstream_waitrequest;
  reg              Medipix_sopc_burst_1_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_1_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_Medipix_sopc_burst_1_downstream_latency_counter;
  wire             pre_flush_Medipix_sopc_burst_1_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module) & (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module) & ((~Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_1_downstream_read | (1 & ~d1_cpu_linux_jtag_debug_module_end_xfer & Medipix_sopc_burst_1_downstream_read))) & ((~Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module | ~Medipix_sopc_burst_1_downstream_write | (1 & Medipix_sopc_burst_1_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_1_downstream_address_to_slave = Medipix_sopc_burst_1_downstream_address;

  //Medipix_sopc_burst_1_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_read_but_no_slave_selected <= 0;
      else 
        Medipix_sopc_burst_1_downstream_read_but_no_slave_selected <= Medipix_sopc_burst_1_downstream_read & Medipix_sopc_burst_1_downstream_run & ~Medipix_sopc_burst_1_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign Medipix_sopc_burst_1_downstream_is_granted_some_slave = Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_1_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_1_downstream_readdatavalid = Medipix_sopc_burst_1_downstream_read_but_no_slave_selected |
    pre_flush_Medipix_sopc_burst_1_downstream_readdatavalid |
    Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module;

  //Medipix_sopc_burst_1/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_1_downstream_readdata = cpu_linux_jtag_debug_module_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_waitrequest = ~Medipix_sopc_burst_1_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_latency_counter <= 0;
      else 
        Medipix_sopc_burst_1_downstream_latency_counter <= p1_Medipix_sopc_burst_1_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_Medipix_sopc_burst_1_downstream_latency_counter = ((Medipix_sopc_burst_1_downstream_run & Medipix_sopc_burst_1_downstream_read))? latency_load_value :
    (Medipix_sopc_burst_1_downstream_latency_counter)? Medipix_sopc_burst_1_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //Medipix_sopc_burst_1_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_1_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_1_downstream_address_last_time <= Medipix_sopc_burst_1_downstream_address;
    end


  //Medipix_sopc_burst_1/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_1_downstream_waitrequest & (Medipix_sopc_burst_1_downstream_read | Medipix_sopc_burst_1_downstream_write);
    end


  //Medipix_sopc_burst_1_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_1_downstream_address != Medipix_sopc_burst_1_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_1_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_1_downstream_burstcount_last_time <= Medipix_sopc_burst_1_downstream_burstcount;
    end


  //Medipix_sopc_burst_1_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_1_downstream_burstcount != Medipix_sopc_burst_1_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_1_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_1_downstream_byteenable_last_time <= Medipix_sopc_burst_1_downstream_byteenable;
    end


  //Medipix_sopc_burst_1_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_1_downstream_byteenable != Medipix_sopc_burst_1_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_1_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_1_downstream_read_last_time <= Medipix_sopc_burst_1_downstream_read;
    end


  //Medipix_sopc_burst_1_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_1_downstream_read != Medipix_sopc_burst_1_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_1_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_1_downstream_write_last_time <= Medipix_sopc_burst_1_downstream_write;
    end


  //Medipix_sopc_burst_1_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_1_downstream_write != Medipix_sopc_burst_1_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_1_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_1_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_1_downstream_writedata_last_time <= Medipix_sopc_burst_1_downstream_writedata;
    end


  //Medipix_sopc_burst_1_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_1_downstream_writedata != Medipix_sopc_burst_1_downstream_writedata_last_time) & Medipix_sopc_burst_1_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_1_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_10_upstream_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_10_upstream_module (
                                                                                     // inputs:
                                                                                      clear_fifo,
                                                                                      clk,
                                                                                      data_in,
                                                                                      read,
                                                                                      reset_n,
                                                                                      sync_reset,
                                                                                      write,

                                                                                     // outputs:
                                                                                      data_out,
                                                                                      empty,
                                                                                      fifo_contains_ones_n,
                                                                                      full
                                                                                   )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_10_upstream_arbitrator (
                                                   // inputs:
                                                    Medipix_sopc_burst_10_upstream_readdata,
                                                    Medipix_sopc_burst_10_upstream_readdatavalid,
                                                    Medipix_sopc_burst_10_upstream_waitrequest,
                                                    clk,
                                                    cpu_linux_data_master_address_to_slave,
                                                    cpu_linux_data_master_burstcount,
                                                    cpu_linux_data_master_byteenable,
                                                    cpu_linux_data_master_debugaccess,
                                                    cpu_linux_data_master_latency_counter,
                                                    cpu_linux_data_master_read,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                    cpu_linux_data_master_write,
                                                    cpu_linux_data_master_writedata,
                                                    reset_n,

                                                   // outputs:
                                                    Medipix_sopc_burst_10_upstream_address,
                                                    Medipix_sopc_burst_10_upstream_burstcount,
                                                    Medipix_sopc_burst_10_upstream_byteaddress,
                                                    Medipix_sopc_burst_10_upstream_byteenable,
                                                    Medipix_sopc_burst_10_upstream_debugaccess,
                                                    Medipix_sopc_burst_10_upstream_read,
                                                    Medipix_sopc_burst_10_upstream_readdata_from_sa,
                                                    Medipix_sopc_burst_10_upstream_waitrequest_from_sa,
                                                    Medipix_sopc_burst_10_upstream_write,
                                                    Medipix_sopc_burst_10_upstream_writedata,
                                                    cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream,
                                                    cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                    cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream,
                                                    d1_Medipix_sopc_burst_10_upstream_end_xfer
                                                 )
;

  output  [  3: 0] Medipix_sopc_burst_10_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_10_upstream_burstcount;
  output  [  4: 0] Medipix_sopc_burst_10_upstream_byteaddress;
  output  [  1: 0] Medipix_sopc_burst_10_upstream_byteenable;
  output           Medipix_sopc_burst_10_upstream_debugaccess;
  output           Medipix_sopc_burst_10_upstream_read;
  output  [ 15: 0] Medipix_sopc_burst_10_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_10_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_10_upstream_write;
  output  [ 15: 0] Medipix_sopc_burst_10_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream;
  output           d1_Medipix_sopc_burst_10_upstream_end_xfer;
  input   [ 15: 0] Medipix_sopc_burst_10_upstream_readdata;
  input            Medipix_sopc_burst_10_upstream_readdatavalid;
  input            Medipix_sopc_burst_10_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [  3: 0] Medipix_sopc_burst_10_upstream_address;
  wire             Medipix_sopc_burst_10_upstream_allgrants;
  wire             Medipix_sopc_burst_10_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_10_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_10_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_10_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_10_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_10_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_10_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_10_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_burstcount;
  wire             Medipix_sopc_burst_10_upstream_burstcount_fifo_empty;
  wire    [  4: 0] Medipix_sopc_burst_10_upstream_byteaddress;
  wire    [  1: 0] Medipix_sopc_burst_10_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_10_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_10_upstream_debugaccess;
  wire             Medipix_sopc_burst_10_upstream_end_xfer;
  wire             Medipix_sopc_burst_10_upstream_firsttransfer;
  wire             Medipix_sopc_burst_10_upstream_grant_vector;
  wire             Medipix_sopc_burst_10_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_10_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_10_upstream_load_fifo;
  wire             Medipix_sopc_burst_10_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_10_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_10_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_next_burst_count;
  wire             Medipix_sopc_burst_10_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_10_upstream_read;
  wire    [ 15: 0] Medipix_sopc_burst_10_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_10_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_10_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_10_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_10_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_10_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_10_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_10_upstream_waits_for_read;
  wire             Medipix_sopc_burst_10_upstream_waits_for_write;
  wire             Medipix_sopc_burst_10_upstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_10_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_10_upstream;
  reg              d1_Medipix_sopc_burst_10_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_10_upstream_load_fifo;
  wire    [ 27: 0] shifted_address_to_Medipix_sopc_burst_10_upstream_from_cpu_linux_data_master;
  wire             wait_for_Medipix_sopc_burst_10_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_10_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_10_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream));
  //assign Medipix_sopc_burst_10_upstream_readdatavalid_from_sa = Medipix_sopc_burst_10_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_readdatavalid_from_sa = Medipix_sopc_burst_10_upstream_readdatavalid;

  //assign Medipix_sopc_burst_10_upstream_readdata_from_sa = Medipix_sopc_burst_10_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_readdata_from_sa = Medipix_sopc_burst_10_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream = ({cpu_linux_data_master_address_to_slave[27 : 5] , 5'b0} == 28'h8000040) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_10_upstream_waitrequest_from_sa = Medipix_sopc_burst_10_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_waitrequest_from_sa = Medipix_sopc_burst_10_upstream_waitrequest;

  //Medipix_sopc_burst_10_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_10_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_10_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_10_upstream;

  //Medipix_sopc_burst_10_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_arb_share_counter_next_value = Medipix_sopc_burst_10_upstream_firsttransfer ? (Medipix_sopc_burst_10_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_10_upstream_arb_share_counter ? (Medipix_sopc_burst_10_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_10_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_allgrants = |Medipix_sopc_burst_10_upstream_grant_vector;

  //Medipix_sopc_burst_10_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_end_xfer = ~(Medipix_sopc_burst_10_upstream_waits_for_read | Medipix_sopc_burst_10_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream = Medipix_sopc_burst_10_upstream_end_xfer & (~Medipix_sopc_burst_10_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_10_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream & Medipix_sopc_burst_10_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream & ~Medipix_sopc_burst_10_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_10_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_10_upstream_arb_counter_enable)
          Medipix_sopc_burst_10_upstream_arb_share_counter <= Medipix_sopc_burst_10_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_10_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_10_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_10_upstream & ~Medipix_sopc_burst_10_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_10_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_10_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_10/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_10_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_10_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_10_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_10/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_10_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_10_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_10_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_move_on_to_next_transaction = Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_10_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_10_upstream, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_10_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_10_upstream_module burstcount_fifo_for_Medipix_sopc_burst_10_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_10_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_10_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_10_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read & Medipix_sopc_burst_10_upstream_load_fifo & ~(Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_10_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_10_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_current_burst_minus_one = Medipix_sopc_burst_10_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_10_upstream, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read) & ~Medipix_sopc_burst_10_upstream_load_fifo))? Medipix_sopc_burst_10_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read & Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_10_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_10_upstream_selected_burstcount :
    (Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_10_upstream_transaction_burst_count :
    Medipix_sopc_burst_10_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_10_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_10_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_10_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read)))
          Medipix_sopc_burst_10_upstream_current_burst <= Medipix_sopc_burst_10_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_10_upstream_load_fifo = (~Medipix_sopc_burst_10_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read) & Medipix_sopc_burst_10_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_10_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read) & ~Medipix_sopc_burst_10_upstream_load_fifo | Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_10_upstream_load_fifo <= p0_Medipix_sopc_burst_10_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_10_upstream, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_10_upstream_current_burst_minus_one) & Medipix_sopc_burst_10_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_10_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_10_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_10_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_10_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_10_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_10_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_10_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_10_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream = Medipix_sopc_burst_10_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_10_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_10/upstream, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_10/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_10_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream;

  //allow new arb cycle for Medipix_sopc_burst_10/upstream, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_10_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_10_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_10_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_firsttransfer = Medipix_sopc_burst_10_upstream_begins_xfer ? Medipix_sopc_burst_10_upstream_unreg_firsttransfer : Medipix_sopc_burst_10_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_10_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_10_upstream_slavearbiterlockenable & Medipix_sopc_burst_10_upstream_any_continuerequest);

  //Medipix_sopc_burst_10_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_10_upstream_begins_xfer)
          Medipix_sopc_burst_10_upstream_reg_firsttransfer <= Medipix_sopc_burst_10_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_10_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_10_upstream_write) && (Medipix_sopc_burst_10_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_10_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_10_upstream_read) && (Medipix_sopc_burst_10_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_10_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_10_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_10_upstream_begins_xfer)
          Medipix_sopc_burst_10_upstream_bbt_burstcounter <= Medipix_sopc_burst_10_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_10_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_beginbursttransfer_internal = Medipix_sopc_burst_10_upstream_begins_xfer & (Medipix_sopc_burst_10_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_10_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_10_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream & cpu_linux_data_master_write;

  assign shifted_address_to_Medipix_sopc_burst_10_upstream_from_cpu_linux_data_master = cpu_linux_data_master_address_to_slave;
  //Medipix_sopc_burst_10_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_address = shifted_address_to_Medipix_sopc_burst_10_upstream_from_cpu_linux_data_master >> 2;

  //d1_Medipix_sopc_burst_10_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_10_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_10_upstream_end_xfer <= Medipix_sopc_burst_10_upstream_end_xfer;
    end


  //Medipix_sopc_burst_10_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_waits_for_read = Medipix_sopc_burst_10_upstream_in_a_read_cycle & Medipix_sopc_burst_10_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_10_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_10_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_10_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_waits_for_write = Medipix_sopc_burst_10_upstream_in_a_write_cycle & Medipix_sopc_burst_10_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_10_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_10_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_10_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_10_upstream_counter = 0;
  //Medipix_sopc_burst_10_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_10_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_10/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_10/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_10_downstream_arbitrator (
                                                     // inputs:
                                                      Medipix_sopc_burst_10_downstream_address,
                                                      Medipix_sopc_burst_10_downstream_burstcount,
                                                      Medipix_sopc_burst_10_downstream_byteenable,
                                                      Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port,
                                                      Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port,
                                                      Medipix_sopc_burst_10_downstream_read,
                                                      Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port,
                                                      Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port,
                                                      Medipix_sopc_burst_10_downstream_write,
                                                      Medipix_sopc_burst_10_downstream_writedata,
                                                      clk,
                                                      d1_spi_0_spi_control_port_end_xfer,
                                                      reset_n,
                                                      spi_0_spi_control_port_readdata_from_sa,

                                                     // outputs:
                                                      Medipix_sopc_burst_10_downstream_address_to_slave,
                                                      Medipix_sopc_burst_10_downstream_latency_counter,
                                                      Medipix_sopc_burst_10_downstream_readdata,
                                                      Medipix_sopc_burst_10_downstream_readdatavalid,
                                                      Medipix_sopc_burst_10_downstream_reset_n,
                                                      Medipix_sopc_burst_10_downstream_waitrequest
                                                   )
;

  output  [  3: 0] Medipix_sopc_burst_10_downstream_address_to_slave;
  output           Medipix_sopc_burst_10_downstream_latency_counter;
  output  [ 15: 0] Medipix_sopc_burst_10_downstream_readdata;
  output           Medipix_sopc_burst_10_downstream_readdatavalid;
  output           Medipix_sopc_burst_10_downstream_reset_n;
  output           Medipix_sopc_burst_10_downstream_waitrequest;
  input   [  3: 0] Medipix_sopc_burst_10_downstream_address;
  input            Medipix_sopc_burst_10_downstream_burstcount;
  input   [  1: 0] Medipix_sopc_burst_10_downstream_byteenable;
  input            Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port;
  input            Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port;
  input            Medipix_sopc_burst_10_downstream_read;
  input            Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port;
  input            Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port;
  input            Medipix_sopc_burst_10_downstream_write;
  input   [ 15: 0] Medipix_sopc_burst_10_downstream_writedata;
  input            clk;
  input            d1_spi_0_spi_control_port_end_xfer;
  input            reset_n;
  input   [ 15: 0] spi_0_spi_control_port_readdata_from_sa;

  reg     [  3: 0] Medipix_sopc_burst_10_downstream_address_last_time;
  wire    [  3: 0] Medipix_sopc_burst_10_downstream_address_to_slave;
  reg              Medipix_sopc_burst_10_downstream_burstcount_last_time;
  reg     [  1: 0] Medipix_sopc_burst_10_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_10_downstream_latency_counter;
  reg              Medipix_sopc_burst_10_downstream_read_last_time;
  wire    [ 15: 0] Medipix_sopc_burst_10_downstream_readdata;
  wire             Medipix_sopc_burst_10_downstream_readdatavalid;
  wire             Medipix_sopc_burst_10_downstream_reset_n;
  wire             Medipix_sopc_burst_10_downstream_run;
  wire             Medipix_sopc_burst_10_downstream_waitrequest;
  reg              Medipix_sopc_burst_10_downstream_write_last_time;
  reg     [ 15: 0] Medipix_sopc_burst_10_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             pre_flush_Medipix_sopc_burst_10_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port | ~Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port) & ((~Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port | ~(Medipix_sopc_burst_10_downstream_read | Medipix_sopc_burst_10_downstream_write) | (1 & ~d1_spi_0_spi_control_port_end_xfer & (Medipix_sopc_burst_10_downstream_read | Medipix_sopc_burst_10_downstream_write)))) & ((~Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port | ~(Medipix_sopc_burst_10_downstream_read | Medipix_sopc_burst_10_downstream_write) | (1 & ~d1_spi_0_spi_control_port_end_xfer & (Medipix_sopc_burst_10_downstream_read | Medipix_sopc_burst_10_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_10_downstream_address_to_slave = Medipix_sopc_burst_10_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_10_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_10_downstream_readdatavalid = 0 |
    pre_flush_Medipix_sopc_burst_10_downstream_readdatavalid |
    Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port;

  //Medipix_sopc_burst_10/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_10_downstream_readdata = spi_0_spi_control_port_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_waitrequest = ~Medipix_sopc_burst_10_downstream_run;

  //latent max counter, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_latency_counter = 0;

  //Medipix_sopc_burst_10_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_10_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_10_downstream_address_last_time <= Medipix_sopc_burst_10_downstream_address;
    end


  //Medipix_sopc_burst_10/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_10_downstream_waitrequest & (Medipix_sopc_burst_10_downstream_read | Medipix_sopc_burst_10_downstream_write);
    end


  //Medipix_sopc_burst_10_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_10_downstream_address != Medipix_sopc_burst_10_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_10_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_10_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_10_downstream_burstcount_last_time <= Medipix_sopc_burst_10_downstream_burstcount;
    end


  //Medipix_sopc_burst_10_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_10_downstream_burstcount != Medipix_sopc_burst_10_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_10_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_10_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_10_downstream_byteenable_last_time <= Medipix_sopc_burst_10_downstream_byteenable;
    end


  //Medipix_sopc_burst_10_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_10_downstream_byteenable != Medipix_sopc_burst_10_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_10_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_10_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_10_downstream_read_last_time <= Medipix_sopc_burst_10_downstream_read;
    end


  //Medipix_sopc_burst_10_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_10_downstream_read != Medipix_sopc_burst_10_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_10_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_10_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_10_downstream_write_last_time <= Medipix_sopc_burst_10_downstream_write;
    end


  //Medipix_sopc_burst_10_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_10_downstream_write != Medipix_sopc_burst_10_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_10_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_10_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_10_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_10_downstream_writedata_last_time <= Medipix_sopc_burst_10_downstream_writedata;
    end


  //Medipix_sopc_burst_10_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_10_downstream_writedata != Medipix_sopc_burst_10_downstream_writedata_last_time) & Medipix_sopc_burst_10_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_10_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_11_upstream_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_11_upstream_module (
                                                                                     // inputs:
                                                                                      clear_fifo,
                                                                                      clk,
                                                                                      data_in,
                                                                                      read,
                                                                                      reset_n,
                                                                                      sync_reset,
                                                                                      write,

                                                                                     // outputs:
                                                                                      data_out,
                                                                                      empty,
                                                                                      fifo_contains_ones_n,
                                                                                      full
                                                                                   )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_11_upstream_arbitrator (
                                                   // inputs:
                                                    Medipix_sopc_burst_11_upstream_readdata,
                                                    Medipix_sopc_burst_11_upstream_readdatavalid,
                                                    Medipix_sopc_burst_11_upstream_waitrequest,
                                                    clk,
                                                    cpu_linux_data_master_address_to_slave,
                                                    cpu_linux_data_master_burstcount,
                                                    cpu_linux_data_master_byteenable,
                                                    cpu_linux_data_master_debugaccess,
                                                    cpu_linux_data_master_latency_counter,
                                                    cpu_linux_data_master_read,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                    cpu_linux_data_master_write,
                                                    cpu_linux_data_master_writedata,
                                                    reset_n,

                                                   // outputs:
                                                    Medipix_sopc_burst_11_upstream_address,
                                                    Medipix_sopc_burst_11_upstream_burstcount,
                                                    Medipix_sopc_burst_11_upstream_byteaddress,
                                                    Medipix_sopc_burst_11_upstream_byteenable,
                                                    Medipix_sopc_burst_11_upstream_debugaccess,
                                                    Medipix_sopc_burst_11_upstream_read,
                                                    Medipix_sopc_burst_11_upstream_readdata_from_sa,
                                                    Medipix_sopc_burst_11_upstream_waitrequest_from_sa,
                                                    Medipix_sopc_burst_11_upstream_write,
                                                    Medipix_sopc_burst_11_upstream_writedata,
                                                    cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream,
                                                    cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream,
                                                    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                    cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream,
                                                    d1_Medipix_sopc_burst_11_upstream_end_xfer
                                                 )
;

  output  [  3: 0] Medipix_sopc_burst_11_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_11_upstream_burstcount;
  output  [  4: 0] Medipix_sopc_burst_11_upstream_byteaddress;
  output  [  1: 0] Medipix_sopc_burst_11_upstream_byteenable;
  output           Medipix_sopc_burst_11_upstream_debugaccess;
  output           Medipix_sopc_burst_11_upstream_read;
  output  [ 15: 0] Medipix_sopc_burst_11_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_11_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_11_upstream_write;
  output  [ 15: 0] Medipix_sopc_burst_11_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream;
  output           d1_Medipix_sopc_burst_11_upstream_end_xfer;
  input   [ 15: 0] Medipix_sopc_burst_11_upstream_readdata;
  input            Medipix_sopc_burst_11_upstream_readdatavalid;
  input            Medipix_sopc_burst_11_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [  3: 0] Medipix_sopc_burst_11_upstream_address;
  wire             Medipix_sopc_burst_11_upstream_allgrants;
  wire             Medipix_sopc_burst_11_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_11_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_11_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_11_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_11_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_11_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_11_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_11_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_burstcount;
  wire             Medipix_sopc_burst_11_upstream_burstcount_fifo_empty;
  wire    [  4: 0] Medipix_sopc_burst_11_upstream_byteaddress;
  wire    [  1: 0] Medipix_sopc_burst_11_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_11_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_11_upstream_debugaccess;
  wire             Medipix_sopc_burst_11_upstream_end_xfer;
  wire             Medipix_sopc_burst_11_upstream_firsttransfer;
  wire             Medipix_sopc_burst_11_upstream_grant_vector;
  wire             Medipix_sopc_burst_11_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_11_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_11_upstream_load_fifo;
  wire             Medipix_sopc_burst_11_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_11_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_11_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_next_burst_count;
  wire             Medipix_sopc_burst_11_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_11_upstream_read;
  wire    [ 15: 0] Medipix_sopc_burst_11_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_11_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_11_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_11_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_11_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_11_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_11_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_11_upstream_waits_for_read;
  wire             Medipix_sopc_burst_11_upstream_waits_for_write;
  wire             Medipix_sopc_burst_11_upstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_11_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_11_upstream;
  reg              d1_Medipix_sopc_burst_11_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_11_upstream_load_fifo;
  wire    [ 27: 0] shifted_address_to_Medipix_sopc_burst_11_upstream_from_cpu_linux_data_master;
  wire             wait_for_Medipix_sopc_burst_11_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_11_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_11_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream));
  //assign Medipix_sopc_burst_11_upstream_readdatavalid_from_sa = Medipix_sopc_burst_11_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_readdatavalid_from_sa = Medipix_sopc_burst_11_upstream_readdatavalid;

  //assign Medipix_sopc_burst_11_upstream_readdata_from_sa = Medipix_sopc_burst_11_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_readdata_from_sa = Medipix_sopc_burst_11_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream = ({cpu_linux_data_master_address_to_slave[27 : 5] , 5'b0} == 28'h8000020) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_11_upstream_waitrequest_from_sa = Medipix_sopc_burst_11_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_waitrequest_from_sa = Medipix_sopc_burst_11_upstream_waitrequest;

  //Medipix_sopc_burst_11_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_11_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_11_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_11_upstream;

  //Medipix_sopc_burst_11_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_arb_share_counter_next_value = Medipix_sopc_burst_11_upstream_firsttransfer ? (Medipix_sopc_burst_11_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_11_upstream_arb_share_counter ? (Medipix_sopc_burst_11_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_11_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_allgrants = |Medipix_sopc_burst_11_upstream_grant_vector;

  //Medipix_sopc_burst_11_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_end_xfer = ~(Medipix_sopc_burst_11_upstream_waits_for_read | Medipix_sopc_burst_11_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream = Medipix_sopc_burst_11_upstream_end_xfer & (~Medipix_sopc_burst_11_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_11_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream & Medipix_sopc_burst_11_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream & ~Medipix_sopc_burst_11_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_11_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_11_upstream_arb_counter_enable)
          Medipix_sopc_burst_11_upstream_arb_share_counter <= Medipix_sopc_burst_11_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_11_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_11_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_11_upstream & ~Medipix_sopc_burst_11_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_11_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_11_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_11/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_11_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_11_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_11_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_11/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_11_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_11_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_11_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_move_on_to_next_transaction = Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_11_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_11_upstream, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_11_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_11_upstream_module burstcount_fifo_for_Medipix_sopc_burst_11_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_11_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_11_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_11_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read & Medipix_sopc_burst_11_upstream_load_fifo & ~(Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_11_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_11_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_current_burst_minus_one = Medipix_sopc_burst_11_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_11_upstream, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read) & ~Medipix_sopc_burst_11_upstream_load_fifo))? Medipix_sopc_burst_11_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read & Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_11_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_11_upstream_selected_burstcount :
    (Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_11_upstream_transaction_burst_count :
    Medipix_sopc_burst_11_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_11_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_11_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_11_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read)))
          Medipix_sopc_burst_11_upstream_current_burst <= Medipix_sopc_burst_11_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_11_upstream_load_fifo = (~Medipix_sopc_burst_11_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read) & Medipix_sopc_burst_11_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_11_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read) & ~Medipix_sopc_burst_11_upstream_load_fifo | Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_11_upstream_load_fifo <= p0_Medipix_sopc_burst_11_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_11_upstream, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_11_upstream_current_burst_minus_one) & Medipix_sopc_burst_11_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_11_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_11_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_11_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_11_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_11_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_11_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_11_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_11_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream = Medipix_sopc_burst_11_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_11_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_11/upstream, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_11/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_11_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream;

  //allow new arb cycle for Medipix_sopc_burst_11/upstream, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_11_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_11_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_11_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_firsttransfer = Medipix_sopc_burst_11_upstream_begins_xfer ? Medipix_sopc_burst_11_upstream_unreg_firsttransfer : Medipix_sopc_burst_11_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_11_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_11_upstream_slavearbiterlockenable & Medipix_sopc_burst_11_upstream_any_continuerequest);

  //Medipix_sopc_burst_11_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_11_upstream_begins_xfer)
          Medipix_sopc_burst_11_upstream_reg_firsttransfer <= Medipix_sopc_burst_11_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_11_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_11_upstream_write) && (Medipix_sopc_burst_11_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_11_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_11_upstream_read) && (Medipix_sopc_burst_11_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_11_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_11_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_11_upstream_begins_xfer)
          Medipix_sopc_burst_11_upstream_bbt_burstcounter <= Medipix_sopc_burst_11_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_11_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_beginbursttransfer_internal = Medipix_sopc_burst_11_upstream_begins_xfer & (Medipix_sopc_burst_11_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_11_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_11_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream & cpu_linux_data_master_write;

  assign shifted_address_to_Medipix_sopc_burst_11_upstream_from_cpu_linux_data_master = cpu_linux_data_master_address_to_slave;
  //Medipix_sopc_burst_11_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_address = shifted_address_to_Medipix_sopc_burst_11_upstream_from_cpu_linux_data_master >> 2;

  //d1_Medipix_sopc_burst_11_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_11_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_11_upstream_end_xfer <= Medipix_sopc_burst_11_upstream_end_xfer;
    end


  //Medipix_sopc_burst_11_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_waits_for_read = Medipix_sopc_burst_11_upstream_in_a_read_cycle & Medipix_sopc_burst_11_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_11_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_11_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_11_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_waits_for_write = Medipix_sopc_burst_11_upstream_in_a_write_cycle & Medipix_sopc_burst_11_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_11_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_11_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_11_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_11_upstream_counter = 0;
  //Medipix_sopc_burst_11_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_11_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_11/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_11/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_11_downstream_arbitrator (
                                                     // inputs:
                                                      Medipix_sopc_burst_11_downstream_address,
                                                      Medipix_sopc_burst_11_downstream_burstcount,
                                                      Medipix_sopc_burst_11_downstream_byteenable,
                                                      Medipix_sopc_burst_11_downstream_granted_uart_0_s1,
                                                      Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1,
                                                      Medipix_sopc_burst_11_downstream_read,
                                                      Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1,
                                                      Medipix_sopc_burst_11_downstream_requests_uart_0_s1,
                                                      Medipix_sopc_burst_11_downstream_write,
                                                      Medipix_sopc_burst_11_downstream_writedata,
                                                      clk,
                                                      d1_uart_0_s1_end_xfer,
                                                      reset_n,
                                                      uart_0_s1_readdata_from_sa,

                                                     // outputs:
                                                      Medipix_sopc_burst_11_downstream_address_to_slave,
                                                      Medipix_sopc_burst_11_downstream_latency_counter,
                                                      Medipix_sopc_burst_11_downstream_readdata,
                                                      Medipix_sopc_burst_11_downstream_readdatavalid,
                                                      Medipix_sopc_burst_11_downstream_reset_n,
                                                      Medipix_sopc_burst_11_downstream_waitrequest
                                                   )
;

  output  [  3: 0] Medipix_sopc_burst_11_downstream_address_to_slave;
  output           Medipix_sopc_burst_11_downstream_latency_counter;
  output  [ 15: 0] Medipix_sopc_burst_11_downstream_readdata;
  output           Medipix_sopc_burst_11_downstream_readdatavalid;
  output           Medipix_sopc_burst_11_downstream_reset_n;
  output           Medipix_sopc_burst_11_downstream_waitrequest;
  input   [  3: 0] Medipix_sopc_burst_11_downstream_address;
  input            Medipix_sopc_burst_11_downstream_burstcount;
  input   [  1: 0] Medipix_sopc_burst_11_downstream_byteenable;
  input            Medipix_sopc_burst_11_downstream_granted_uart_0_s1;
  input            Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1;
  input            Medipix_sopc_burst_11_downstream_read;
  input            Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1;
  input            Medipix_sopc_burst_11_downstream_requests_uart_0_s1;
  input            Medipix_sopc_burst_11_downstream_write;
  input   [ 15: 0] Medipix_sopc_burst_11_downstream_writedata;
  input            clk;
  input            d1_uart_0_s1_end_xfer;
  input            reset_n;
  input   [ 15: 0] uart_0_s1_readdata_from_sa;

  reg     [  3: 0] Medipix_sopc_burst_11_downstream_address_last_time;
  wire    [  3: 0] Medipix_sopc_burst_11_downstream_address_to_slave;
  reg              Medipix_sopc_burst_11_downstream_burstcount_last_time;
  reg     [  1: 0] Medipix_sopc_burst_11_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_11_downstream_latency_counter;
  reg              Medipix_sopc_burst_11_downstream_read_last_time;
  wire    [ 15: 0] Medipix_sopc_burst_11_downstream_readdata;
  wire             Medipix_sopc_burst_11_downstream_readdatavalid;
  wire             Medipix_sopc_burst_11_downstream_reset_n;
  wire             Medipix_sopc_burst_11_downstream_run;
  wire             Medipix_sopc_burst_11_downstream_waitrequest;
  reg              Medipix_sopc_burst_11_downstream_write_last_time;
  reg     [ 15: 0] Medipix_sopc_burst_11_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             pre_flush_Medipix_sopc_burst_11_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1 | ~Medipix_sopc_burst_11_downstream_requests_uart_0_s1) & ((~Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1 | ~(Medipix_sopc_burst_11_downstream_read | Medipix_sopc_burst_11_downstream_write) | (1 & ~d1_uart_0_s1_end_xfer & (Medipix_sopc_burst_11_downstream_read | Medipix_sopc_burst_11_downstream_write)))) & ((~Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1 | ~(Medipix_sopc_burst_11_downstream_read | Medipix_sopc_burst_11_downstream_write) | (1 & ~d1_uart_0_s1_end_xfer & (Medipix_sopc_burst_11_downstream_read | Medipix_sopc_burst_11_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_11_downstream_address_to_slave = Medipix_sopc_burst_11_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_11_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_11_downstream_readdatavalid = 0 |
    pre_flush_Medipix_sopc_burst_11_downstream_readdatavalid |
    Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1;

  //Medipix_sopc_burst_11/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_11_downstream_readdata = uart_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_waitrequest = ~Medipix_sopc_burst_11_downstream_run;

  //latent max counter, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_latency_counter = 0;

  //Medipix_sopc_burst_11_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_11_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_11_downstream_address_last_time <= Medipix_sopc_burst_11_downstream_address;
    end


  //Medipix_sopc_burst_11/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_11_downstream_waitrequest & (Medipix_sopc_burst_11_downstream_read | Medipix_sopc_burst_11_downstream_write);
    end


  //Medipix_sopc_burst_11_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_11_downstream_address != Medipix_sopc_burst_11_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_11_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_11_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_11_downstream_burstcount_last_time <= Medipix_sopc_burst_11_downstream_burstcount;
    end


  //Medipix_sopc_burst_11_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_11_downstream_burstcount != Medipix_sopc_burst_11_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_11_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_11_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_11_downstream_byteenable_last_time <= Medipix_sopc_burst_11_downstream_byteenable;
    end


  //Medipix_sopc_burst_11_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_11_downstream_byteenable != Medipix_sopc_burst_11_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_11_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_11_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_11_downstream_read_last_time <= Medipix_sopc_burst_11_downstream_read;
    end


  //Medipix_sopc_burst_11_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_11_downstream_read != Medipix_sopc_burst_11_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_11_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_11_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_11_downstream_write_last_time <= Medipix_sopc_burst_11_downstream_write;
    end


  //Medipix_sopc_burst_11_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_11_downstream_write != Medipix_sopc_burst_11_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_11_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_11_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_11_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_11_downstream_writedata_last_time <= Medipix_sopc_burst_11_downstream_writedata;
    end


  //Medipix_sopc_burst_11_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_11_downstream_writedata != Medipix_sopc_burst_11_downstream_writedata_last_time) & Medipix_sopc_burst_11_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_11_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_2_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_2_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_2_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_2_upstream_readdata,
                                                   Medipix_sopc_burst_2_upstream_readdatavalid,
                                                   Medipix_sopc_burst_2_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_2_upstream_address,
                                                   Medipix_sopc_burst_2_upstream_burstcount,
                                                   Medipix_sopc_burst_2_upstream_byteaddress,
                                                   Medipix_sopc_burst_2_upstream_byteenable,
                                                   Medipix_sopc_burst_2_upstream_debugaccess,
                                                   Medipix_sopc_burst_2_upstream_read,
                                                   Medipix_sopc_burst_2_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_2_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_2_upstream_write,
                                                   Medipix_sopc_burst_2_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream,
                                                   d1_Medipix_sopc_burst_2_upstream_end_xfer
                                                )
;

  output  [  2: 0] Medipix_sopc_burst_2_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_2_upstream_burstcount;
  output  [  4: 0] Medipix_sopc_burst_2_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_2_upstream_byteenable;
  output           Medipix_sopc_burst_2_upstream_debugaccess;
  output           Medipix_sopc_burst_2_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_2_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_2_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_2_upstream_write;
  output  [ 31: 0] Medipix_sopc_burst_2_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream;
  output           d1_Medipix_sopc_burst_2_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_2_upstream_readdata;
  input            Medipix_sopc_burst_2_upstream_readdatavalid;
  input            Medipix_sopc_burst_2_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [  2: 0] Medipix_sopc_burst_2_upstream_address;
  wire             Medipix_sopc_burst_2_upstream_allgrants;
  wire             Medipix_sopc_burst_2_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_2_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_2_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_2_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_2_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_2_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_2_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_2_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_burstcount;
  wire             Medipix_sopc_burst_2_upstream_burstcount_fifo_empty;
  wire    [  4: 0] Medipix_sopc_burst_2_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_2_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_2_upstream_debugaccess;
  wire             Medipix_sopc_burst_2_upstream_end_xfer;
  wire             Medipix_sopc_burst_2_upstream_firsttransfer;
  wire             Medipix_sopc_burst_2_upstream_grant_vector;
  wire             Medipix_sopc_burst_2_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_2_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_2_upstream_load_fifo;
  wire             Medipix_sopc_burst_2_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_2_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_2_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_next_burst_count;
  wire             Medipix_sopc_burst_2_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_2_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_2_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_2_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_2_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_2_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_2_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_2_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_2_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_2_upstream_waits_for_read;
  wire             Medipix_sopc_burst_2_upstream_waits_for_write;
  wire             Medipix_sopc_burst_2_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_2_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_2_upstream;
  reg              d1_Medipix_sopc_burst_2_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_2_upstream_load_fifo;
  wire    [ 27: 0] shifted_address_to_Medipix_sopc_burst_2_upstream_from_cpu_linux_data_master;
  wire             wait_for_Medipix_sopc_burst_2_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_2_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_2_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream));
  //assign Medipix_sopc_burst_2_upstream_readdatavalid_from_sa = Medipix_sopc_burst_2_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_readdatavalid_from_sa = Medipix_sopc_burst_2_upstream_readdatavalid;

  //assign Medipix_sopc_burst_2_upstream_readdata_from_sa = Medipix_sopc_burst_2_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_readdata_from_sa = Medipix_sopc_burst_2_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream = ({cpu_linux_data_master_address_to_slave[27 : 3] , 3'b0} == 28'h8001020) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_2_upstream_waitrequest_from_sa = Medipix_sopc_burst_2_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_waitrequest_from_sa = Medipix_sopc_burst_2_upstream_waitrequest;

  //Medipix_sopc_burst_2_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_2_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_2_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_2_upstream;

  //Medipix_sopc_burst_2_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_arb_share_counter_next_value = Medipix_sopc_burst_2_upstream_firsttransfer ? (Medipix_sopc_burst_2_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_2_upstream_arb_share_counter ? (Medipix_sopc_burst_2_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_2_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_allgrants = |Medipix_sopc_burst_2_upstream_grant_vector;

  //Medipix_sopc_burst_2_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_end_xfer = ~(Medipix_sopc_burst_2_upstream_waits_for_read | Medipix_sopc_burst_2_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream = Medipix_sopc_burst_2_upstream_end_xfer & (~Medipix_sopc_burst_2_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_2_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream & Medipix_sopc_burst_2_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream & ~Medipix_sopc_burst_2_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_2_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_2_upstream_arb_counter_enable)
          Medipix_sopc_burst_2_upstream_arb_share_counter <= Medipix_sopc_burst_2_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_2_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_2_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_2_upstream & ~Medipix_sopc_burst_2_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_2_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_2_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_2/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_2_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_2_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_2_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_2/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_2_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_2_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_2_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_move_on_to_next_transaction = Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_2_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_2_upstream, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_2_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_2_upstream_module burstcount_fifo_for_Medipix_sopc_burst_2_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_2_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_2_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_2_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read & Medipix_sopc_burst_2_upstream_load_fifo & ~(Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_2_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_2_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_current_burst_minus_one = Medipix_sopc_burst_2_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_2_upstream, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read) & ~Medipix_sopc_burst_2_upstream_load_fifo))? Medipix_sopc_burst_2_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read & Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_2_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_2_upstream_selected_burstcount :
    (Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_2_upstream_transaction_burst_count :
    Medipix_sopc_burst_2_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_2_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_2_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_2_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read)))
          Medipix_sopc_burst_2_upstream_current_burst <= Medipix_sopc_burst_2_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_2_upstream_load_fifo = (~Medipix_sopc_burst_2_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read) & Medipix_sopc_burst_2_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_2_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read) & ~Medipix_sopc_burst_2_upstream_load_fifo | Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_2_upstream_load_fifo <= p0_Medipix_sopc_burst_2_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_2_upstream, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_2_upstream_current_burst_minus_one) & Medipix_sopc_burst_2_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_2_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_2_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_2_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_2_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_2_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_2_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_2_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_2_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream = Medipix_sopc_burst_2_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_2_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_2/upstream, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_2/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_2_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream;

  //allow new arb cycle for Medipix_sopc_burst_2/upstream, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_2_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_2_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_2_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_firsttransfer = Medipix_sopc_burst_2_upstream_begins_xfer ? Medipix_sopc_burst_2_upstream_unreg_firsttransfer : Medipix_sopc_burst_2_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_2_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_2_upstream_slavearbiterlockenable & Medipix_sopc_burst_2_upstream_any_continuerequest);

  //Medipix_sopc_burst_2_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_2_upstream_begins_xfer)
          Medipix_sopc_burst_2_upstream_reg_firsttransfer <= Medipix_sopc_burst_2_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_2_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_2_upstream_write) && (Medipix_sopc_burst_2_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_2_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_2_upstream_read) && (Medipix_sopc_burst_2_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_2_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_2_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_2_upstream_begins_xfer)
          Medipix_sopc_burst_2_upstream_bbt_burstcounter <= Medipix_sopc_burst_2_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_2_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_beginbursttransfer_internal = Medipix_sopc_burst_2_upstream_begins_xfer & (Medipix_sopc_burst_2_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_2_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_2_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream & cpu_linux_data_master_write;

  assign shifted_address_to_Medipix_sopc_burst_2_upstream_from_cpu_linux_data_master = cpu_linux_data_master_address_to_slave;
  //Medipix_sopc_burst_2_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_address = shifted_address_to_Medipix_sopc_burst_2_upstream_from_cpu_linux_data_master >> 2;

  //d1_Medipix_sopc_burst_2_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_2_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_2_upstream_end_xfer <= Medipix_sopc_burst_2_upstream_end_xfer;
    end


  //Medipix_sopc_burst_2_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_waits_for_read = Medipix_sopc_burst_2_upstream_in_a_read_cycle & Medipix_sopc_burst_2_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_2_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_2_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_2_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_waits_for_write = Medipix_sopc_burst_2_upstream_in_a_write_cycle & Medipix_sopc_burst_2_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_2_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_2_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_2_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_2_upstream_counter = 0;
  //Medipix_sopc_burst_2_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_2_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_2/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_2/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_2_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_2_downstream_address,
                                                     Medipix_sopc_burst_2_downstream_burstcount,
                                                     Medipix_sopc_burst_2_downstream_byteenable,
                                                     Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave,
                                                     Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave,
                                                     Medipix_sopc_burst_2_downstream_read,
                                                     Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave,
                                                     Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave,
                                                     Medipix_sopc_burst_2_downstream_write,
                                                     Medipix_sopc_burst_2_downstream_writedata,
                                                     clk,
                                                     d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
                                                     jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
                                                     jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_2_downstream_address_to_slave,
                                                     Medipix_sopc_burst_2_downstream_latency_counter,
                                                     Medipix_sopc_burst_2_downstream_readdata,
                                                     Medipix_sopc_burst_2_downstream_readdatavalid,
                                                     Medipix_sopc_burst_2_downstream_reset_n,
                                                     Medipix_sopc_burst_2_downstream_waitrequest
                                                  )
;

  output  [  2: 0] Medipix_sopc_burst_2_downstream_address_to_slave;
  output           Medipix_sopc_burst_2_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_2_downstream_readdata;
  output           Medipix_sopc_burst_2_downstream_readdatavalid;
  output           Medipix_sopc_burst_2_downstream_reset_n;
  output           Medipix_sopc_burst_2_downstream_waitrequest;
  input   [  2: 0] Medipix_sopc_burst_2_downstream_address;
  input            Medipix_sopc_burst_2_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_2_downstream_byteenable;
  input            Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave;
  input            Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave;
  input            Medipix_sopc_burst_2_downstream_read;
  input            Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  input            Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave;
  input            Medipix_sopc_burst_2_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_2_downstream_writedata;
  input            clk;
  input            d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  input   [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  input            reset_n;

  reg     [  2: 0] Medipix_sopc_burst_2_downstream_address_last_time;
  wire    [  2: 0] Medipix_sopc_burst_2_downstream_address_to_slave;
  reg              Medipix_sopc_burst_2_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_2_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_2_downstream_latency_counter;
  reg              Medipix_sopc_burst_2_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_2_downstream_readdata;
  wire             Medipix_sopc_burst_2_downstream_readdatavalid;
  wire             Medipix_sopc_burst_2_downstream_reset_n;
  wire             Medipix_sopc_burst_2_downstream_run;
  wire             Medipix_sopc_burst_2_downstream_waitrequest;
  reg              Medipix_sopc_burst_2_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_2_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             pre_flush_Medipix_sopc_burst_2_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave | ~Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave) & ((~Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave | ~(Medipix_sopc_burst_2_downstream_read | Medipix_sopc_burst_2_downstream_write) | (1 & ~jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa & (Medipix_sopc_burst_2_downstream_read | Medipix_sopc_burst_2_downstream_write)))) & ((~Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave | ~(Medipix_sopc_burst_2_downstream_read | Medipix_sopc_burst_2_downstream_write) | (1 & ~jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa & (Medipix_sopc_burst_2_downstream_read | Medipix_sopc_burst_2_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_2_downstream_address_to_slave = Medipix_sopc_burst_2_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_2_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_2_downstream_readdatavalid = 0 |
    pre_flush_Medipix_sopc_burst_2_downstream_readdatavalid |
    Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave;

  //Medipix_sopc_burst_2/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_2_downstream_readdata = jtag_uart_0_avalon_jtag_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_waitrequest = ~Medipix_sopc_burst_2_downstream_run;

  //latent max counter, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_latency_counter = 0;

  //Medipix_sopc_burst_2_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_2_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_2_downstream_address_last_time <= Medipix_sopc_burst_2_downstream_address;
    end


  //Medipix_sopc_burst_2/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_2_downstream_waitrequest & (Medipix_sopc_burst_2_downstream_read | Medipix_sopc_burst_2_downstream_write);
    end


  //Medipix_sopc_burst_2_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_2_downstream_address != Medipix_sopc_burst_2_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_2_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_2_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_2_downstream_burstcount_last_time <= Medipix_sopc_burst_2_downstream_burstcount;
    end


  //Medipix_sopc_burst_2_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_2_downstream_burstcount != Medipix_sopc_burst_2_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_2_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_2_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_2_downstream_byteenable_last_time <= Medipix_sopc_burst_2_downstream_byteenable;
    end


  //Medipix_sopc_burst_2_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_2_downstream_byteenable != Medipix_sopc_burst_2_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_2_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_2_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_2_downstream_read_last_time <= Medipix_sopc_burst_2_downstream_read;
    end


  //Medipix_sopc_burst_2_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_2_downstream_read != Medipix_sopc_burst_2_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_2_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_2_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_2_downstream_write_last_time <= Medipix_sopc_burst_2_downstream_write;
    end


  //Medipix_sopc_burst_2_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_2_downstream_write != Medipix_sopc_burst_2_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_2_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_2_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_2_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_2_downstream_writedata_last_time <= Medipix_sopc_burst_2_downstream_writedata;
    end


  //Medipix_sopc_burst_2_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_2_downstream_writedata != Medipix_sopc_burst_2_downstream_writedata_last_time) & Medipix_sopc_burst_2_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_2_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_3_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_3_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_3_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_3_upstream_readdata,
                                                   Medipix_sopc_burst_3_upstream_readdatavalid,
                                                   Medipix_sopc_burst_3_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_3_upstream_address,
                                                   Medipix_sopc_burst_3_upstream_burstcount,
                                                   Medipix_sopc_burst_3_upstream_byteaddress,
                                                   Medipix_sopc_burst_3_upstream_byteenable,
                                                   Medipix_sopc_burst_3_upstream_debugaccess,
                                                   Medipix_sopc_burst_3_upstream_read,
                                                   Medipix_sopc_burst_3_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_3_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_3_upstream_write,
                                                   Medipix_sopc_burst_3_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream,
                                                   d1_Medipix_sopc_burst_3_upstream_end_xfer
                                                )
;

  output  [  3: 0] Medipix_sopc_burst_3_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_3_upstream_burstcount;
  output  [  4: 0] Medipix_sopc_burst_3_upstream_byteaddress;
  output  [  1: 0] Medipix_sopc_burst_3_upstream_byteenable;
  output           Medipix_sopc_burst_3_upstream_debugaccess;
  output           Medipix_sopc_burst_3_upstream_read;
  output  [ 15: 0] Medipix_sopc_burst_3_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_3_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_3_upstream_write;
  output  [ 15: 0] Medipix_sopc_burst_3_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream;
  output           d1_Medipix_sopc_burst_3_upstream_end_xfer;
  input   [ 15: 0] Medipix_sopc_burst_3_upstream_readdata;
  input            Medipix_sopc_burst_3_upstream_readdatavalid;
  input            Medipix_sopc_burst_3_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [  3: 0] Medipix_sopc_burst_3_upstream_address;
  wire             Medipix_sopc_burst_3_upstream_allgrants;
  wire             Medipix_sopc_burst_3_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_3_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_3_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_3_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_3_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_3_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_3_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_3_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_burstcount;
  wire             Medipix_sopc_burst_3_upstream_burstcount_fifo_empty;
  wire    [  4: 0] Medipix_sopc_burst_3_upstream_byteaddress;
  wire    [  1: 0] Medipix_sopc_burst_3_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_3_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_3_upstream_debugaccess;
  wire             Medipix_sopc_burst_3_upstream_end_xfer;
  wire             Medipix_sopc_burst_3_upstream_firsttransfer;
  wire             Medipix_sopc_burst_3_upstream_grant_vector;
  wire             Medipix_sopc_burst_3_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_3_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_3_upstream_load_fifo;
  wire             Medipix_sopc_burst_3_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_3_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_3_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_next_burst_count;
  wire             Medipix_sopc_burst_3_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_3_upstream_read;
  wire    [ 15: 0] Medipix_sopc_burst_3_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_3_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_3_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_3_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_3_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_3_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_3_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_3_upstream_waits_for_read;
  wire             Medipix_sopc_burst_3_upstream_waits_for_write;
  wire             Medipix_sopc_burst_3_upstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_3_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_3_upstream;
  reg              d1_Medipix_sopc_burst_3_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_3_upstream_load_fifo;
  wire    [ 27: 0] shifted_address_to_Medipix_sopc_burst_3_upstream_from_cpu_linux_data_master;
  wire             wait_for_Medipix_sopc_burst_3_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_3_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_3_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream));
  //assign Medipix_sopc_burst_3_upstream_readdatavalid_from_sa = Medipix_sopc_burst_3_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_readdatavalid_from_sa = Medipix_sopc_burst_3_upstream_readdatavalid;

  //assign Medipix_sopc_burst_3_upstream_readdata_from_sa = Medipix_sopc_burst_3_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_readdata_from_sa = Medipix_sopc_burst_3_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream = ({cpu_linux_data_master_address_to_slave[27 : 5] , 5'b0} == 28'h8001000) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_3_upstream_waitrequest_from_sa = Medipix_sopc_burst_3_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_waitrequest_from_sa = Medipix_sopc_burst_3_upstream_waitrequest;

  //Medipix_sopc_burst_3_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_3_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_3_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_3_upstream;

  //Medipix_sopc_burst_3_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_arb_share_counter_next_value = Medipix_sopc_burst_3_upstream_firsttransfer ? (Medipix_sopc_burst_3_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_3_upstream_arb_share_counter ? (Medipix_sopc_burst_3_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_3_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_allgrants = |Medipix_sopc_burst_3_upstream_grant_vector;

  //Medipix_sopc_burst_3_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_end_xfer = ~(Medipix_sopc_burst_3_upstream_waits_for_read | Medipix_sopc_burst_3_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream = Medipix_sopc_burst_3_upstream_end_xfer & (~Medipix_sopc_burst_3_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_3_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream & Medipix_sopc_burst_3_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream & ~Medipix_sopc_burst_3_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_3_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_3_upstream_arb_counter_enable)
          Medipix_sopc_burst_3_upstream_arb_share_counter <= Medipix_sopc_burst_3_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_3_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_3_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_3_upstream & ~Medipix_sopc_burst_3_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_3_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_3_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_3/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_3_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_3_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_3_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_3/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_3_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_3_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_3_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_move_on_to_next_transaction = Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_3_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_3_upstream, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_3_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_3_upstream_module burstcount_fifo_for_Medipix_sopc_burst_3_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_3_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_3_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_3_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read & Medipix_sopc_burst_3_upstream_load_fifo & ~(Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_3_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_3_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_current_burst_minus_one = Medipix_sopc_burst_3_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_3_upstream, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read) & ~Medipix_sopc_burst_3_upstream_load_fifo))? Medipix_sopc_burst_3_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read & Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_3_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_3_upstream_selected_burstcount :
    (Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_3_upstream_transaction_burst_count :
    Medipix_sopc_burst_3_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_3_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_3_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_3_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read)))
          Medipix_sopc_burst_3_upstream_current_burst <= Medipix_sopc_burst_3_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_3_upstream_load_fifo = (~Medipix_sopc_burst_3_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read) & Medipix_sopc_burst_3_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_3_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read) & ~Medipix_sopc_burst_3_upstream_load_fifo | Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_3_upstream_load_fifo <= p0_Medipix_sopc_burst_3_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_3_upstream, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_3_upstream_current_burst_minus_one) & Medipix_sopc_burst_3_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_3_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_3_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_3_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_3_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_3_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_3_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_3_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_3_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream = Medipix_sopc_burst_3_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_3_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_3/upstream, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_3/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_3_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream;

  //allow new arb cycle for Medipix_sopc_burst_3/upstream, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_3_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_3_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_3_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_firsttransfer = Medipix_sopc_burst_3_upstream_begins_xfer ? Medipix_sopc_burst_3_upstream_unreg_firsttransfer : Medipix_sopc_burst_3_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_3_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_3_upstream_slavearbiterlockenable & Medipix_sopc_burst_3_upstream_any_continuerequest);

  //Medipix_sopc_burst_3_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_3_upstream_begins_xfer)
          Medipix_sopc_burst_3_upstream_reg_firsttransfer <= Medipix_sopc_burst_3_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_3_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_3_upstream_write) && (Medipix_sopc_burst_3_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_3_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_3_upstream_read) && (Medipix_sopc_burst_3_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_3_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_3_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_3_upstream_begins_xfer)
          Medipix_sopc_burst_3_upstream_bbt_burstcounter <= Medipix_sopc_burst_3_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_3_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_beginbursttransfer_internal = Medipix_sopc_burst_3_upstream_begins_xfer & (Medipix_sopc_burst_3_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_3_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_3_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream & cpu_linux_data_master_write;

  assign shifted_address_to_Medipix_sopc_burst_3_upstream_from_cpu_linux_data_master = cpu_linux_data_master_address_to_slave;
  //Medipix_sopc_burst_3_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_address = shifted_address_to_Medipix_sopc_burst_3_upstream_from_cpu_linux_data_master >> 2;

  //d1_Medipix_sopc_burst_3_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_3_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_3_upstream_end_xfer <= Medipix_sopc_burst_3_upstream_end_xfer;
    end


  //Medipix_sopc_burst_3_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_waits_for_read = Medipix_sopc_burst_3_upstream_in_a_read_cycle & Medipix_sopc_burst_3_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_3_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_3_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_3_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_waits_for_write = Medipix_sopc_burst_3_upstream_in_a_write_cycle & Medipix_sopc_burst_3_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_3_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_3_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_3_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_3_upstream_counter = 0;
  //Medipix_sopc_burst_3_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_3_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_3/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_3/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_3_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_3_downstream_address,
                                                     Medipix_sopc_burst_3_downstream_burstcount,
                                                     Medipix_sopc_burst_3_downstream_byteenable,
                                                     Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1,
                                                     Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1,
                                                     Medipix_sopc_burst_3_downstream_read,
                                                     Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1,
                                                     Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1,
                                                     Medipix_sopc_burst_3_downstream_write,
                                                     Medipix_sopc_burst_3_downstream_writedata,
                                                     clk,
                                                     d1_sys_clk_freq_s1_end_xfer,
                                                     reset_n,
                                                     sys_clk_freq_s1_readdata_from_sa,

                                                    // outputs:
                                                     Medipix_sopc_burst_3_downstream_address_to_slave,
                                                     Medipix_sopc_burst_3_downstream_latency_counter,
                                                     Medipix_sopc_burst_3_downstream_readdata,
                                                     Medipix_sopc_burst_3_downstream_readdatavalid,
                                                     Medipix_sopc_burst_3_downstream_reset_n,
                                                     Medipix_sopc_burst_3_downstream_waitrequest
                                                  )
;

  output  [  3: 0] Medipix_sopc_burst_3_downstream_address_to_slave;
  output           Medipix_sopc_burst_3_downstream_latency_counter;
  output  [ 15: 0] Medipix_sopc_burst_3_downstream_readdata;
  output           Medipix_sopc_burst_3_downstream_readdatavalid;
  output           Medipix_sopc_burst_3_downstream_reset_n;
  output           Medipix_sopc_burst_3_downstream_waitrequest;
  input   [  3: 0] Medipix_sopc_burst_3_downstream_address;
  input            Medipix_sopc_burst_3_downstream_burstcount;
  input   [  1: 0] Medipix_sopc_burst_3_downstream_byteenable;
  input            Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1;
  input            Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1;
  input            Medipix_sopc_burst_3_downstream_read;
  input            Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1;
  input            Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1;
  input            Medipix_sopc_burst_3_downstream_write;
  input   [ 15: 0] Medipix_sopc_burst_3_downstream_writedata;
  input            clk;
  input            d1_sys_clk_freq_s1_end_xfer;
  input            reset_n;
  input   [ 15: 0] sys_clk_freq_s1_readdata_from_sa;

  reg     [  3: 0] Medipix_sopc_burst_3_downstream_address_last_time;
  wire    [  3: 0] Medipix_sopc_burst_3_downstream_address_to_slave;
  reg              Medipix_sopc_burst_3_downstream_burstcount_last_time;
  reg     [  1: 0] Medipix_sopc_burst_3_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_3_downstream_latency_counter;
  reg              Medipix_sopc_burst_3_downstream_read_last_time;
  wire    [ 15: 0] Medipix_sopc_burst_3_downstream_readdata;
  wire             Medipix_sopc_burst_3_downstream_readdatavalid;
  wire             Medipix_sopc_burst_3_downstream_reset_n;
  wire             Medipix_sopc_burst_3_downstream_run;
  wire             Medipix_sopc_burst_3_downstream_waitrequest;
  reg              Medipix_sopc_burst_3_downstream_write_last_time;
  reg     [ 15: 0] Medipix_sopc_burst_3_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             pre_flush_Medipix_sopc_burst_3_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1 | ~Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1) & ((~Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1 | ~Medipix_sopc_burst_3_downstream_read | (1 & ~d1_sys_clk_freq_s1_end_xfer & Medipix_sopc_burst_3_downstream_read))) & ((~Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1 | ~Medipix_sopc_burst_3_downstream_write | (1 & Medipix_sopc_burst_3_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_3_downstream_address_to_slave = Medipix_sopc_burst_3_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_3_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_3_downstream_readdatavalid = 0 |
    pre_flush_Medipix_sopc_burst_3_downstream_readdatavalid |
    Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1;

  //Medipix_sopc_burst_3/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_3_downstream_readdata = sys_clk_freq_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_waitrequest = ~Medipix_sopc_burst_3_downstream_run;

  //latent max counter, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_latency_counter = 0;

  //Medipix_sopc_burst_3_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_3_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_3_downstream_address_last_time <= Medipix_sopc_burst_3_downstream_address;
    end


  //Medipix_sopc_burst_3/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_3_downstream_waitrequest & (Medipix_sopc_burst_3_downstream_read | Medipix_sopc_burst_3_downstream_write);
    end


  //Medipix_sopc_burst_3_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_3_downstream_address != Medipix_sopc_burst_3_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_3_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_3_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_3_downstream_burstcount_last_time <= Medipix_sopc_burst_3_downstream_burstcount;
    end


  //Medipix_sopc_burst_3_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_3_downstream_burstcount != Medipix_sopc_burst_3_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_3_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_3_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_3_downstream_byteenable_last_time <= Medipix_sopc_burst_3_downstream_byteenable;
    end


  //Medipix_sopc_burst_3_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_3_downstream_byteenable != Medipix_sopc_burst_3_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_3_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_3_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_3_downstream_read_last_time <= Medipix_sopc_burst_3_downstream_read;
    end


  //Medipix_sopc_burst_3_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_3_downstream_read != Medipix_sopc_burst_3_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_3_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_3_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_3_downstream_write_last_time <= Medipix_sopc_burst_3_downstream_write;
    end


  //Medipix_sopc_burst_3_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_3_downstream_write != Medipix_sopc_burst_3_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_3_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_3_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_3_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_3_downstream_writedata_last_time <= Medipix_sopc_burst_3_downstream_writedata;
    end


  //Medipix_sopc_burst_3_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_3_downstream_writedata != Medipix_sopc_burst_3_downstream_writedata_last_time) & Medipix_sopc_burst_3_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_3_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_4_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  3: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  3: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  3: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  3: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  3: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  3: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  3: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  3: 0] p17_stage_17;
  wire             p18_full_18;
  wire    [  3: 0] p18_stage_18;
  wire             p19_full_19;
  wire    [  3: 0] p19_stage_19;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p20_full_20;
  wire    [  3: 0] p20_stage_20;
  wire             p21_full_21;
  wire    [  3: 0] p21_stage_21;
  wire             p22_full_22;
  wire    [  3: 0] p22_stage_22;
  wire             p23_full_23;
  wire    [  3: 0] p23_stage_23;
  wire             p24_full_24;
  wire    [  3: 0] p24_stage_24;
  wire             p25_full_25;
  wire    [  3: 0] p25_stage_25;
  wire             p26_full_26;
  wire    [  3: 0] p26_stage_26;
  wire             p27_full_27;
  wire    [  3: 0] p27_stage_27;
  wire             p28_full_28;
  wire    [  3: 0] p28_stage_28;
  wire             p29_full_29;
  wire    [  3: 0] p29_stage_29;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p30_full_30;
  wire    [  3: 0] p30_stage_30;
  wire             p31_full_31;
  wire    [  3: 0] p31_stage_31;
  wire             p32_full_32;
  wire    [  3: 0] p32_stage_32;
  wire             p33_full_33;
  wire    [  3: 0] p33_stage_33;
  wire             p34_full_34;
  wire    [  3: 0] p34_stage_34;
  wire             p35_full_35;
  wire    [  3: 0] p35_stage_35;
  wire             p36_full_36;
  wire    [  3: 0] p36_stage_36;
  wire             p37_full_37;
  wire    [  3: 0] p37_stage_37;
  wire             p38_full_38;
  wire    [  3: 0] p38_stage_38;
  wire             p39_full_39;
  wire    [  3: 0] p39_stage_39;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p40_full_40;
  wire    [  3: 0] p40_stage_40;
  wire             p41_full_41;
  wire    [  3: 0] p41_stage_41;
  wire             p42_full_42;
  wire    [  3: 0] p42_stage_42;
  wire             p43_full_43;
  wire    [  3: 0] p43_stage_43;
  wire             p44_full_44;
  wire    [  3: 0] p44_stage_44;
  wire             p45_full_45;
  wire    [  3: 0] p45_stage_45;
  wire             p46_full_46;
  wire    [  3: 0] p46_stage_46;
  wire             p47_full_47;
  wire    [  3: 0] p47_stage_47;
  wire             p48_full_48;
  wire    [  3: 0] p48_stage_48;
  wire             p49_full_49;
  wire    [  3: 0] p49_stage_49;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p50_full_50;
  wire    [  3: 0] p50_stage_50;
  wire             p51_full_51;
  wire    [  3: 0] p51_stage_51;
  wire             p52_full_52;
  wire    [  3: 0] p52_stage_52;
  wire             p53_full_53;
  wire    [  3: 0] p53_stage_53;
  wire             p54_full_54;
  wire    [  3: 0] p54_stage_54;
  wire             p55_full_55;
  wire    [  3: 0] p55_stage_55;
  wire             p56_full_56;
  wire    [  3: 0] p56_stage_56;
  wire             p57_full_57;
  wire    [  3: 0] p57_stage_57;
  wire             p58_full_58;
  wire    [  3: 0] p58_stage_58;
  wire             p59_full_59;
  wire    [  3: 0] p59_stage_59;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p60_full_60;
  wire    [  3: 0] p60_stage_60;
  wire             p61_full_61;
  wire    [  3: 0] p61_stage_61;
  wire             p62_full_62;
  wire    [  3: 0] p62_stage_62;
  wire             p63_full_63;
  wire    [  3: 0] p63_stage_63;
  wire             p64_full_64;
  wire    [  3: 0] p64_stage_64;
  wire             p65_full_65;
  wire    [  3: 0] p65_stage_65;
  wire             p66_full_66;
  wire    [  3: 0] p66_stage_66;
  wire             p67_full_67;
  wire    [  3: 0] p67_stage_67;
  wire             p68_full_68;
  wire    [  3: 0] p68_stage_68;
  wire             p69_full_69;
  wire    [  3: 0] p69_stage_69;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p70_full_70;
  wire    [  3: 0] p70_stage_70;
  wire             p71_full_71;
  wire    [  3: 0] p71_stage_71;
  wire             p72_full_72;
  wire    [  3: 0] p72_stage_72;
  wire             p73_full_73;
  wire    [  3: 0] p73_stage_73;
  wire             p74_full_74;
  wire    [  3: 0] p74_stage_74;
  wire             p75_full_75;
  wire    [  3: 0] p75_stage_75;
  wire             p76_full_76;
  wire    [  3: 0] p76_stage_76;
  wire             p77_full_77;
  wire    [  3: 0] p77_stage_77;
  wire             p78_full_78;
  wire    [  3: 0] p78_stage_78;
  wire             p79_full_79;
  wire    [  3: 0] p79_stage_79;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p80_full_80;
  wire    [  3: 0] p80_stage_80;
  wire             p81_full_81;
  wire    [  3: 0] p81_stage_81;
  wire             p82_full_82;
  wire    [  3: 0] p82_stage_82;
  wire             p83_full_83;
  wire    [  3: 0] p83_stage_83;
  wire             p84_full_84;
  wire    [  3: 0] p84_stage_84;
  wire             p85_full_85;
  wire    [  3: 0] p85_stage_85;
  wire             p86_full_86;
  wire    [  3: 0] p86_stage_86;
  wire             p87_full_87;
  wire    [  3: 0] p87_stage_87;
  wire             p88_full_88;
  wire    [  3: 0] p88_stage_88;
  wire             p89_full_89;
  wire    [  3: 0] p89_stage_89;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  wire             p90_full_90;
  wire    [  3: 0] p90_stage_90;
  wire             p91_full_91;
  wire    [  3: 0] p91_stage_91;
  wire             p92_full_92;
  wire    [  3: 0] p92_stage_92;
  wire             p93_full_93;
  wire    [  3: 0] p93_stage_93;
  wire             p94_full_94;
  wire    [  3: 0] p94_stage_94;
  wire             p95_full_95;
  wire    [  3: 0] p95_stage_95;
  wire             p96_full_96;
  wire    [  3: 0] p96_stage_96;
  wire             p97_full_97;
  wire    [  3: 0] p97_stage_97;
  wire             p9_full_9;
  wire    [  3: 0] p9_stage_9;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_10;
  reg     [  3: 0] stage_11;
  reg     [  3: 0] stage_12;
  reg     [  3: 0] stage_13;
  reg     [  3: 0] stage_14;
  reg     [  3: 0] stage_15;
  reg     [  3: 0] stage_16;
  reg     [  3: 0] stage_17;
  reg     [  3: 0] stage_18;
  reg     [  3: 0] stage_19;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_20;
  reg     [  3: 0] stage_21;
  reg     [  3: 0] stage_22;
  reg     [  3: 0] stage_23;
  reg     [  3: 0] stage_24;
  reg     [  3: 0] stage_25;
  reg     [  3: 0] stage_26;
  reg     [  3: 0] stage_27;
  reg     [  3: 0] stage_28;
  reg     [  3: 0] stage_29;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_30;
  reg     [  3: 0] stage_31;
  reg     [  3: 0] stage_32;
  reg     [  3: 0] stage_33;
  reg     [  3: 0] stage_34;
  reg     [  3: 0] stage_35;
  reg     [  3: 0] stage_36;
  reg     [  3: 0] stage_37;
  reg     [  3: 0] stage_38;
  reg     [  3: 0] stage_39;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_40;
  reg     [  3: 0] stage_41;
  reg     [  3: 0] stage_42;
  reg     [  3: 0] stage_43;
  reg     [  3: 0] stage_44;
  reg     [  3: 0] stage_45;
  reg     [  3: 0] stage_46;
  reg     [  3: 0] stage_47;
  reg     [  3: 0] stage_48;
  reg     [  3: 0] stage_49;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_50;
  reg     [  3: 0] stage_51;
  reg     [  3: 0] stage_52;
  reg     [  3: 0] stage_53;
  reg     [  3: 0] stage_54;
  reg     [  3: 0] stage_55;
  reg     [  3: 0] stage_56;
  reg     [  3: 0] stage_57;
  reg     [  3: 0] stage_58;
  reg     [  3: 0] stage_59;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_60;
  reg     [  3: 0] stage_61;
  reg     [  3: 0] stage_62;
  reg     [  3: 0] stage_63;
  reg     [  3: 0] stage_64;
  reg     [  3: 0] stage_65;
  reg     [  3: 0] stage_66;
  reg     [  3: 0] stage_67;
  reg     [  3: 0] stage_68;
  reg     [  3: 0] stage_69;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_70;
  reg     [  3: 0] stage_71;
  reg     [  3: 0] stage_72;
  reg     [  3: 0] stage_73;
  reg     [  3: 0] stage_74;
  reg     [  3: 0] stage_75;
  reg     [  3: 0] stage_76;
  reg     [  3: 0] stage_77;
  reg     [  3: 0] stage_78;
  reg     [  3: 0] stage_79;
  reg     [  3: 0] stage_8;
  reg     [  3: 0] stage_80;
  reg     [  3: 0] stage_81;
  reg     [  3: 0] stage_82;
  reg     [  3: 0] stage_83;
  reg     [  3: 0] stage_84;
  reg     [  3: 0] stage_85;
  reg     [  3: 0] stage_86;
  reg     [  3: 0] stage_87;
  reg     [  3: 0] stage_88;
  reg     [  3: 0] stage_89;
  reg     [  3: 0] stage_9;
  reg     [  3: 0] stage_90;
  reg     [  3: 0] stage_91;
  reg     [  3: 0] stage_92;
  reg     [  3: 0] stage_93;
  reg     [  3: 0] stage_94;
  reg     [  3: 0] stage_95;
  reg     [  3: 0] stage_96;
  reg     [  3: 0] stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_4_upstream_module (
                                                                                           // inputs:
                                                                                            clear_fifo,
                                                                                            clk,
                                                                                            data_in,
                                                                                            read,
                                                                                            reset_n,
                                                                                            sync_reset,
                                                                                            write,

                                                                                           // outputs:
                                                                                            data_out,
                                                                                            empty,
                                                                                            fifo_contains_ones_n,
                                                                                            full
                                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p96_full_96;
  wire             p96_stage_96;
  wire             p97_full_97;
  wire             p97_stage_97;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  reg              stage_96;
  reg              stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_4_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_4_upstream_readdata,
                                                   Medipix_sopc_burst_4_upstream_readdatavalid,
                                                   Medipix_sopc_burst_4_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_instruction_master_address_to_slave,
                                                   cpu_linux_instruction_master_burstcount,
                                                   cpu_linux_instruction_master_latency_counter,
                                                   cpu_linux_instruction_master_read,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_4_upstream_address,
                                                   Medipix_sopc_burst_4_upstream_byteaddress,
                                                   Medipix_sopc_burst_4_upstream_byteenable,
                                                   Medipix_sopc_burst_4_upstream_debugaccess,
                                                   Medipix_sopc_burst_4_upstream_read,
                                                   Medipix_sopc_burst_4_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_4_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_4_upstream_write,
                                                   cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream,
                                                   cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register,
                                                   cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream,
                                                   d1_Medipix_sopc_burst_4_upstream_end_xfer
                                                )
;

  output  [ 26: 0] Medipix_sopc_burst_4_upstream_address;
  output  [ 28: 0] Medipix_sopc_burst_4_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_4_upstream_byteenable;
  output           Medipix_sopc_burst_4_upstream_debugaccess;
  output           Medipix_sopc_burst_4_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_4_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_4_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_4_upstream_write;
  output           cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream;
  output           cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream;
  output           cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream;
  output           cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register;
  output           cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream;
  output           d1_Medipix_sopc_burst_4_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_4_upstream_readdata;
  input            Medipix_sopc_burst_4_upstream_readdatavalid;
  input            Medipix_sopc_burst_4_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_instruction_master_address_to_slave;
  input   [  3: 0] cpu_linux_instruction_master_burstcount;
  input            cpu_linux_instruction_master_latency_counter;
  input            cpu_linux_instruction_master_read;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register;
  input            reset_n;

  wire    [ 26: 0] Medipix_sopc_burst_4_upstream_address;
  wire             Medipix_sopc_burst_4_upstream_allgrants;
  wire             Medipix_sopc_burst_4_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_4_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_4_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_4_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_4_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_arb_share_set_values;
  wire             Medipix_sopc_burst_4_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_4_upstream_begins_xfer;
  wire             Medipix_sopc_burst_4_upstream_burstcount_fifo_empty;
  wire    [ 28: 0] Medipix_sopc_burst_4_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_4_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_4_upstream_debugaccess;
  wire             Medipix_sopc_burst_4_upstream_end_xfer;
  wire             Medipix_sopc_burst_4_upstream_firsttransfer;
  wire             Medipix_sopc_burst_4_upstream_grant_vector;
  wire             Medipix_sopc_burst_4_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_4_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_4_upstream_load_fifo;
  wire             Medipix_sopc_burst_4_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_4_upstream_move_on_to_next_transaction;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_next_burst_count;
  wire             Medipix_sopc_burst_4_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_4_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_4_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_4_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_4_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_4_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_4_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_4_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_4_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_4_upstream_waits_for_read;
  wire             Medipix_sopc_burst_4_upstream_waits_for_write;
  wire             Medipix_sopc_burst_4_upstream_write;
  wire             cpu_linux_instruction_master_arbiterlock;
  wire             cpu_linux_instruction_master_arbiterlock2;
  wire             cpu_linux_instruction_master_continuerequest;
  wire             cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_rdv_fifo_output_from_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register;
  wire             cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_4_upstream;
  reg              d1_Medipix_sopc_burst_4_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_4_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_4_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_4_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_4_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream));
  //assign Medipix_sopc_burst_4_upstream_readdatavalid_from_sa = Medipix_sopc_burst_4_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_readdatavalid_from_sa = Medipix_sopc_burst_4_upstream_readdatavalid;

  //assign Medipix_sopc_burst_4_upstream_readdata_from_sa = Medipix_sopc_burst_4_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_readdata_from_sa = Medipix_sopc_burst_4_upstream_readdata;

  assign cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream = (({cpu_linux_instruction_master_address_to_slave[27] , 27'b0} == 28'h0) & (cpu_linux_instruction_master_read)) & cpu_linux_instruction_master_read;
  //assign Medipix_sopc_burst_4_upstream_waitrequest_from_sa = Medipix_sopc_burst_4_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_waitrequest_from_sa = Medipix_sopc_burst_4_upstream_waitrequest;

  //Medipix_sopc_burst_4_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_arb_share_set_values = 1;

  //Medipix_sopc_burst_4_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_4_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_any_bursting_master_saved_grant = cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_4_upstream;

  //Medipix_sopc_burst_4_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_arb_share_counter_next_value = Medipix_sopc_burst_4_upstream_firsttransfer ? (Medipix_sopc_burst_4_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_4_upstream_arb_share_counter ? (Medipix_sopc_burst_4_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_4_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_allgrants = |Medipix_sopc_burst_4_upstream_grant_vector;

  //Medipix_sopc_burst_4_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_end_xfer = ~(Medipix_sopc_burst_4_upstream_waits_for_read | Medipix_sopc_burst_4_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream = Medipix_sopc_burst_4_upstream_end_xfer & (~Medipix_sopc_burst_4_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_4_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream & Medipix_sopc_burst_4_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream & ~Medipix_sopc_burst_4_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_4_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_4_upstream_arb_counter_enable)
          Medipix_sopc_burst_4_upstream_arb_share_counter <= Medipix_sopc_burst_4_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_4_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_4_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_4_upstream & ~Medipix_sopc_burst_4_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_4_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_4_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/instruction_master Medipix_sopc_burst_4/upstream arbiterlock, which is an e_assign
  assign cpu_linux_instruction_master_arbiterlock = Medipix_sopc_burst_4_upstream_slavearbiterlockenable & cpu_linux_instruction_master_continuerequest;

  //Medipix_sopc_burst_4_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_4_upstream_arb_share_counter_next_value;

  //cpu_linux/instruction_master Medipix_sopc_burst_4/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_instruction_master_arbiterlock2 = Medipix_sopc_burst_4_upstream_slavearbiterlockenable2 & cpu_linux_instruction_master_continuerequest;

  //Medipix_sopc_burst_4_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_any_continuerequest = 1;

  //cpu_linux_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_instruction_master_continuerequest = 1;

  assign cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream = cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream & ~((cpu_linux_instruction_master_read & ((cpu_linux_instruction_master_latency_counter != 0) | (1 < cpu_linux_instruction_master_latency_counter) | (|cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register) | (|cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_4_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_move_on_to_next_transaction = Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_4_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_4_upstream, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_selected_burstcount = (cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream)? cpu_linux_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_4_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_4_upstream_module burstcount_fifo_for_Medipix_sopc_burst_4_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_4_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_4_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_4_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read & Medipix_sopc_burst_4_upstream_load_fifo & ~(Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_4_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_4_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_current_burst_minus_one = Medipix_sopc_burst_4_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_4_upstream, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read) & ~Medipix_sopc_burst_4_upstream_load_fifo))? Medipix_sopc_burst_4_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read & Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_4_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_4_upstream_selected_burstcount :
    (Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_4_upstream_transaction_burst_count :
    Medipix_sopc_burst_4_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_4_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_4_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_4_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read)))
          Medipix_sopc_burst_4_upstream_current_burst <= Medipix_sopc_burst_4_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_4_upstream_load_fifo = (~Medipix_sopc_burst_4_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read) & Medipix_sopc_burst_4_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_4_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read) & ~Medipix_sopc_burst_4_upstream_load_fifo | Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_4_upstream_load_fifo <= p0_Medipix_sopc_burst_4_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_4_upstream, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_4_upstream_current_burst_minus_one) & Medipix_sopc_burst_4_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_4_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_4_upstream_module rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_4_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream),
      .data_out             (cpu_linux_instruction_master_rdv_fifo_output_from_Medipix_sopc_burst_4_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_4_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_4_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_4_upstream_waits_for_read)
    );

  assign cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register = ~cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_4_upstream;
  //local readdatavalid cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream, which is an e_mux
  assign cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream = Medipix_sopc_burst_4_upstream_readdatavalid_from_sa;

  //byteaddress mux for Medipix_sopc_burst_4/upstream, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_byteaddress = cpu_linux_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream = cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream;

  //cpu_linux/instruction_master saved-grant Medipix_sopc_burst_4/upstream, which is an e_assign
  assign cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_4_upstream = cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream;

  //allow new arb cycle for Medipix_sopc_burst_4/upstream, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_4_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_4_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_4_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_firsttransfer = Medipix_sopc_burst_4_upstream_begins_xfer ? Medipix_sopc_burst_4_upstream_unreg_firsttransfer : Medipix_sopc_burst_4_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_4_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_4_upstream_slavearbiterlockenable & Medipix_sopc_burst_4_upstream_any_continuerequest);

  //Medipix_sopc_burst_4_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_4_upstream_begins_xfer)
          Medipix_sopc_burst_4_upstream_reg_firsttransfer <= Medipix_sopc_burst_4_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_4_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_beginbursttransfer_internal = Medipix_sopc_burst_4_upstream_begins_xfer;

  //Medipix_sopc_burst_4_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_read = cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream & cpu_linux_instruction_master_read;

  //Medipix_sopc_burst_4_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_write = 0;

  //Medipix_sopc_burst_4_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_address = cpu_linux_instruction_master_address_to_slave;

  //d1_Medipix_sopc_burst_4_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_4_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_4_upstream_end_xfer <= Medipix_sopc_burst_4_upstream_end_xfer;
    end


  //Medipix_sopc_burst_4_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_waits_for_read = Medipix_sopc_burst_4_upstream_in_a_read_cycle & Medipix_sopc_burst_4_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_4_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_in_a_read_cycle = cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream & cpu_linux_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_4_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_4_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_waits_for_write = Medipix_sopc_burst_4_upstream_in_a_write_cycle & Medipix_sopc_burst_4_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_4_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_4_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_4_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_4_upstream_counter = 0;
  //Medipix_sopc_burst_4_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_4_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_4/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream && (cpu_linux_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/instruction_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_4/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_4_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_4_downstream_address,
                                                     Medipix_sopc_burst_4_downstream_burstcount,
                                                     Medipix_sopc_burst_4_downstream_byteenable,
                                                     Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1,
                                                     Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1,
                                                     Medipix_sopc_burst_4_downstream_read,
                                                     Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1,
                                                     Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register,
                                                     Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1,
                                                     Medipix_sopc_burst_4_downstream_write,
                                                     Medipix_sopc_burst_4_downstream_writedata,
                                                     clk,
                                                     clock_crossing_s1_readdata_from_sa,
                                                     clock_crossing_s1_waitrequest_from_sa,
                                                     d1_clock_crossing_s1_end_xfer,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_4_downstream_address_to_slave,
                                                     Medipix_sopc_burst_4_downstream_latency_counter,
                                                     Medipix_sopc_burst_4_downstream_readdata,
                                                     Medipix_sopc_burst_4_downstream_readdatavalid,
                                                     Medipix_sopc_burst_4_downstream_reset_n,
                                                     Medipix_sopc_burst_4_downstream_waitrequest
                                                  )
;

  output  [ 26: 0] Medipix_sopc_burst_4_downstream_address_to_slave;
  output           Medipix_sopc_burst_4_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_4_downstream_readdata;
  output           Medipix_sopc_burst_4_downstream_readdatavalid;
  output           Medipix_sopc_burst_4_downstream_reset_n;
  output           Medipix_sopc_burst_4_downstream_waitrequest;
  input   [ 26: 0] Medipix_sopc_burst_4_downstream_address;
  input            Medipix_sopc_burst_4_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_4_downstream_byteenable;
  input            Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1;
  input            Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1;
  input            Medipix_sopc_burst_4_downstream_read;
  input            Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1;
  input            Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register;
  input            Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1;
  input            Medipix_sopc_burst_4_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_4_downstream_writedata;
  input            clk;
  input   [ 31: 0] clock_crossing_s1_readdata_from_sa;
  input            clock_crossing_s1_waitrequest_from_sa;
  input            d1_clock_crossing_s1_end_xfer;
  input            reset_n;

  reg     [ 26: 0] Medipix_sopc_burst_4_downstream_address_last_time;
  wire    [ 26: 0] Medipix_sopc_burst_4_downstream_address_to_slave;
  reg              Medipix_sopc_burst_4_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_4_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_4_downstream_is_granted_some_slave;
  reg              Medipix_sopc_burst_4_downstream_latency_counter;
  reg              Medipix_sopc_burst_4_downstream_read_but_no_slave_selected;
  reg              Medipix_sopc_burst_4_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_4_downstream_readdata;
  wire             Medipix_sopc_burst_4_downstream_readdatavalid;
  wire             Medipix_sopc_burst_4_downstream_reset_n;
  wire             Medipix_sopc_burst_4_downstream_run;
  wire             Medipix_sopc_burst_4_downstream_waitrequest;
  reg              Medipix_sopc_burst_4_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_4_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_Medipix_sopc_burst_4_downstream_latency_counter;
  wire             pre_flush_Medipix_sopc_burst_4_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1 | ~Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1) & (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 | ~Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1) & ((~Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1 | ~(Medipix_sopc_burst_4_downstream_read | Medipix_sopc_burst_4_downstream_write) | (1 & ~clock_crossing_s1_waitrequest_from_sa & (Medipix_sopc_burst_4_downstream_read | Medipix_sopc_burst_4_downstream_write)))) & ((~Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1 | ~(Medipix_sopc_burst_4_downstream_read | Medipix_sopc_burst_4_downstream_write) | (1 & ~clock_crossing_s1_waitrequest_from_sa & (Medipix_sopc_burst_4_downstream_read | Medipix_sopc_burst_4_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_4_downstream_address_to_slave = Medipix_sopc_burst_4_downstream_address;

  //Medipix_sopc_burst_4_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_read_but_no_slave_selected <= 0;
      else 
        Medipix_sopc_burst_4_downstream_read_but_no_slave_selected <= Medipix_sopc_burst_4_downstream_read & Medipix_sopc_burst_4_downstream_run & ~Medipix_sopc_burst_4_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign Medipix_sopc_burst_4_downstream_is_granted_some_slave = Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_4_downstream_readdatavalid = Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_4_downstream_readdatavalid = Medipix_sopc_burst_4_downstream_read_but_no_slave_selected |
    pre_flush_Medipix_sopc_burst_4_downstream_readdatavalid;

  //Medipix_sopc_burst_4/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_4_downstream_readdata = clock_crossing_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_waitrequest = ~Medipix_sopc_burst_4_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_latency_counter <= 0;
      else 
        Medipix_sopc_burst_4_downstream_latency_counter <= p1_Medipix_sopc_burst_4_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_Medipix_sopc_burst_4_downstream_latency_counter = ((Medipix_sopc_burst_4_downstream_run & Medipix_sopc_burst_4_downstream_read))? latency_load_value :
    (Medipix_sopc_burst_4_downstream_latency_counter)? Medipix_sopc_burst_4_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //Medipix_sopc_burst_4_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_4_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_4_downstream_address_last_time <= Medipix_sopc_burst_4_downstream_address;
    end


  //Medipix_sopc_burst_4/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_4_downstream_waitrequest & (Medipix_sopc_burst_4_downstream_read | Medipix_sopc_burst_4_downstream_write);
    end


  //Medipix_sopc_burst_4_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_4_downstream_address != Medipix_sopc_burst_4_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_4_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_4_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_4_downstream_burstcount_last_time <= Medipix_sopc_burst_4_downstream_burstcount;
    end


  //Medipix_sopc_burst_4_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_4_downstream_burstcount != Medipix_sopc_burst_4_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_4_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_4_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_4_downstream_byteenable_last_time <= Medipix_sopc_burst_4_downstream_byteenable;
    end


  //Medipix_sopc_burst_4_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_4_downstream_byteenable != Medipix_sopc_burst_4_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_4_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_4_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_4_downstream_read_last_time <= Medipix_sopc_burst_4_downstream_read;
    end


  //Medipix_sopc_burst_4_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_4_downstream_read != Medipix_sopc_burst_4_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_4_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_4_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_4_downstream_write_last_time <= Medipix_sopc_burst_4_downstream_write;
    end


  //Medipix_sopc_burst_4_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_4_downstream_write != Medipix_sopc_burst_4_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_4_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_4_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_4_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_4_downstream_writedata_last_time <= Medipix_sopc_burst_4_downstream_writedata;
    end


  //Medipix_sopc_burst_4_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_4_downstream_writedata != Medipix_sopc_burst_4_downstream_writedata_last_time) & Medipix_sopc_burst_4_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_4_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_5_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  3: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  3: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  3: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  3: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  3: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  3: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  3: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  3: 0] p17_stage_17;
  wire             p18_full_18;
  wire    [  3: 0] p18_stage_18;
  wire             p19_full_19;
  wire    [  3: 0] p19_stage_19;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p20_full_20;
  wire    [  3: 0] p20_stage_20;
  wire             p21_full_21;
  wire    [  3: 0] p21_stage_21;
  wire             p22_full_22;
  wire    [  3: 0] p22_stage_22;
  wire             p23_full_23;
  wire    [  3: 0] p23_stage_23;
  wire             p24_full_24;
  wire    [  3: 0] p24_stage_24;
  wire             p25_full_25;
  wire    [  3: 0] p25_stage_25;
  wire             p26_full_26;
  wire    [  3: 0] p26_stage_26;
  wire             p27_full_27;
  wire    [  3: 0] p27_stage_27;
  wire             p28_full_28;
  wire    [  3: 0] p28_stage_28;
  wire             p29_full_29;
  wire    [  3: 0] p29_stage_29;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p30_full_30;
  wire    [  3: 0] p30_stage_30;
  wire             p31_full_31;
  wire    [  3: 0] p31_stage_31;
  wire             p32_full_32;
  wire    [  3: 0] p32_stage_32;
  wire             p33_full_33;
  wire    [  3: 0] p33_stage_33;
  wire             p34_full_34;
  wire    [  3: 0] p34_stage_34;
  wire             p35_full_35;
  wire    [  3: 0] p35_stage_35;
  wire             p36_full_36;
  wire    [  3: 0] p36_stage_36;
  wire             p37_full_37;
  wire    [  3: 0] p37_stage_37;
  wire             p38_full_38;
  wire    [  3: 0] p38_stage_38;
  wire             p39_full_39;
  wire    [  3: 0] p39_stage_39;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p40_full_40;
  wire    [  3: 0] p40_stage_40;
  wire             p41_full_41;
  wire    [  3: 0] p41_stage_41;
  wire             p42_full_42;
  wire    [  3: 0] p42_stage_42;
  wire             p43_full_43;
  wire    [  3: 0] p43_stage_43;
  wire             p44_full_44;
  wire    [  3: 0] p44_stage_44;
  wire             p45_full_45;
  wire    [  3: 0] p45_stage_45;
  wire             p46_full_46;
  wire    [  3: 0] p46_stage_46;
  wire             p47_full_47;
  wire    [  3: 0] p47_stage_47;
  wire             p48_full_48;
  wire    [  3: 0] p48_stage_48;
  wire             p49_full_49;
  wire    [  3: 0] p49_stage_49;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p50_full_50;
  wire    [  3: 0] p50_stage_50;
  wire             p51_full_51;
  wire    [  3: 0] p51_stage_51;
  wire             p52_full_52;
  wire    [  3: 0] p52_stage_52;
  wire             p53_full_53;
  wire    [  3: 0] p53_stage_53;
  wire             p54_full_54;
  wire    [  3: 0] p54_stage_54;
  wire             p55_full_55;
  wire    [  3: 0] p55_stage_55;
  wire             p56_full_56;
  wire    [  3: 0] p56_stage_56;
  wire             p57_full_57;
  wire    [  3: 0] p57_stage_57;
  wire             p58_full_58;
  wire    [  3: 0] p58_stage_58;
  wire             p59_full_59;
  wire    [  3: 0] p59_stage_59;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p60_full_60;
  wire    [  3: 0] p60_stage_60;
  wire             p61_full_61;
  wire    [  3: 0] p61_stage_61;
  wire             p62_full_62;
  wire    [  3: 0] p62_stage_62;
  wire             p63_full_63;
  wire    [  3: 0] p63_stage_63;
  wire             p64_full_64;
  wire    [  3: 0] p64_stage_64;
  wire             p65_full_65;
  wire    [  3: 0] p65_stage_65;
  wire             p66_full_66;
  wire    [  3: 0] p66_stage_66;
  wire             p67_full_67;
  wire    [  3: 0] p67_stage_67;
  wire             p68_full_68;
  wire    [  3: 0] p68_stage_68;
  wire             p69_full_69;
  wire    [  3: 0] p69_stage_69;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p70_full_70;
  wire    [  3: 0] p70_stage_70;
  wire             p71_full_71;
  wire    [  3: 0] p71_stage_71;
  wire             p72_full_72;
  wire    [  3: 0] p72_stage_72;
  wire             p73_full_73;
  wire    [  3: 0] p73_stage_73;
  wire             p74_full_74;
  wire    [  3: 0] p74_stage_74;
  wire             p75_full_75;
  wire    [  3: 0] p75_stage_75;
  wire             p76_full_76;
  wire    [  3: 0] p76_stage_76;
  wire             p77_full_77;
  wire    [  3: 0] p77_stage_77;
  wire             p78_full_78;
  wire    [  3: 0] p78_stage_78;
  wire             p79_full_79;
  wire    [  3: 0] p79_stage_79;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p80_full_80;
  wire    [  3: 0] p80_stage_80;
  wire             p81_full_81;
  wire    [  3: 0] p81_stage_81;
  wire             p82_full_82;
  wire    [  3: 0] p82_stage_82;
  wire             p83_full_83;
  wire    [  3: 0] p83_stage_83;
  wire             p84_full_84;
  wire    [  3: 0] p84_stage_84;
  wire             p85_full_85;
  wire    [  3: 0] p85_stage_85;
  wire             p86_full_86;
  wire    [  3: 0] p86_stage_86;
  wire             p87_full_87;
  wire    [  3: 0] p87_stage_87;
  wire             p88_full_88;
  wire    [  3: 0] p88_stage_88;
  wire             p89_full_89;
  wire    [  3: 0] p89_stage_89;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  wire             p90_full_90;
  wire    [  3: 0] p90_stage_90;
  wire             p91_full_91;
  wire    [  3: 0] p91_stage_91;
  wire             p92_full_92;
  wire    [  3: 0] p92_stage_92;
  wire             p93_full_93;
  wire    [  3: 0] p93_stage_93;
  wire             p94_full_94;
  wire    [  3: 0] p94_stage_94;
  wire             p95_full_95;
  wire    [  3: 0] p95_stage_95;
  wire             p96_full_96;
  wire    [  3: 0] p96_stage_96;
  wire             p97_full_97;
  wire    [  3: 0] p97_stage_97;
  wire             p9_full_9;
  wire    [  3: 0] p9_stage_9;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_10;
  reg     [  3: 0] stage_11;
  reg     [  3: 0] stage_12;
  reg     [  3: 0] stage_13;
  reg     [  3: 0] stage_14;
  reg     [  3: 0] stage_15;
  reg     [  3: 0] stage_16;
  reg     [  3: 0] stage_17;
  reg     [  3: 0] stage_18;
  reg     [  3: 0] stage_19;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_20;
  reg     [  3: 0] stage_21;
  reg     [  3: 0] stage_22;
  reg     [  3: 0] stage_23;
  reg     [  3: 0] stage_24;
  reg     [  3: 0] stage_25;
  reg     [  3: 0] stage_26;
  reg     [  3: 0] stage_27;
  reg     [  3: 0] stage_28;
  reg     [  3: 0] stage_29;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_30;
  reg     [  3: 0] stage_31;
  reg     [  3: 0] stage_32;
  reg     [  3: 0] stage_33;
  reg     [  3: 0] stage_34;
  reg     [  3: 0] stage_35;
  reg     [  3: 0] stage_36;
  reg     [  3: 0] stage_37;
  reg     [  3: 0] stage_38;
  reg     [  3: 0] stage_39;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_40;
  reg     [  3: 0] stage_41;
  reg     [  3: 0] stage_42;
  reg     [  3: 0] stage_43;
  reg     [  3: 0] stage_44;
  reg     [  3: 0] stage_45;
  reg     [  3: 0] stage_46;
  reg     [  3: 0] stage_47;
  reg     [  3: 0] stage_48;
  reg     [  3: 0] stage_49;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_50;
  reg     [  3: 0] stage_51;
  reg     [  3: 0] stage_52;
  reg     [  3: 0] stage_53;
  reg     [  3: 0] stage_54;
  reg     [  3: 0] stage_55;
  reg     [  3: 0] stage_56;
  reg     [  3: 0] stage_57;
  reg     [  3: 0] stage_58;
  reg     [  3: 0] stage_59;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_60;
  reg     [  3: 0] stage_61;
  reg     [  3: 0] stage_62;
  reg     [  3: 0] stage_63;
  reg     [  3: 0] stage_64;
  reg     [  3: 0] stage_65;
  reg     [  3: 0] stage_66;
  reg     [  3: 0] stage_67;
  reg     [  3: 0] stage_68;
  reg     [  3: 0] stage_69;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_70;
  reg     [  3: 0] stage_71;
  reg     [  3: 0] stage_72;
  reg     [  3: 0] stage_73;
  reg     [  3: 0] stage_74;
  reg     [  3: 0] stage_75;
  reg     [  3: 0] stage_76;
  reg     [  3: 0] stage_77;
  reg     [  3: 0] stage_78;
  reg     [  3: 0] stage_79;
  reg     [  3: 0] stage_8;
  reg     [  3: 0] stage_80;
  reg     [  3: 0] stage_81;
  reg     [  3: 0] stage_82;
  reg     [  3: 0] stage_83;
  reg     [  3: 0] stage_84;
  reg     [  3: 0] stage_85;
  reg     [  3: 0] stage_86;
  reg     [  3: 0] stage_87;
  reg     [  3: 0] stage_88;
  reg     [  3: 0] stage_89;
  reg     [  3: 0] stage_9;
  reg     [  3: 0] stage_90;
  reg     [  3: 0] stage_91;
  reg     [  3: 0] stage_92;
  reg     [  3: 0] stage_93;
  reg     [  3: 0] stage_94;
  reg     [  3: 0] stage_95;
  reg     [  3: 0] stage_96;
  reg     [  3: 0] stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_5_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  reg              full_96;
  reg              full_97;
  wire             full_98;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p96_full_96;
  wire             p96_stage_96;
  wire             p97_full_97;
  wire             p97_stage_97;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  reg              stage_96;
  reg              stage_97;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_97;
  assign empty = !full_0;
  assign full_98 = 0;
  //data_97, which is an e_mux
  assign p97_stage_97 = ((full_98 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_97 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_97))
          if (sync_reset & full_97 & !((full_98 == 0) & read & write))
              stage_97 <= 0;
          else 
            stage_97 <= p97_stage_97;
    end


  //control_97, which is an e_mux
  assign p97_full_97 = ((read & !write) == 0)? full_96 :
    0;

  //control_reg_97, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_97 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_97 <= 0;
          else 
            full_97 <= p97_full_97;
    end


  //data_96, which is an e_mux
  assign p96_stage_96 = ((full_97 & ~clear_fifo) == 0)? data_in :
    stage_97;

  //data_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_96 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_96))
          if (sync_reset & full_96 & !((full_97 == 0) & read & write))
              stage_96 <= 0;
          else 
            stage_96 <= p96_stage_96;
    end


  //control_96, which is an e_mux
  assign p96_full_96 = ((read & !write) == 0)? full_95 :
    full_97;

  //control_reg_96, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_96 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_96 <= 0;
          else 
            full_96 <= p96_full_96;
    end


  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    stage_96;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    full_96;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_5_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_5_upstream_readdata,
                                                   Medipix_sopc_burst_5_upstream_readdatavalid,
                                                   Medipix_sopc_burst_5_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_5_upstream_address,
                                                   Medipix_sopc_burst_5_upstream_burstcount,
                                                   Medipix_sopc_burst_5_upstream_byteaddress,
                                                   Medipix_sopc_burst_5_upstream_byteenable,
                                                   Medipix_sopc_burst_5_upstream_debugaccess,
                                                   Medipix_sopc_burst_5_upstream_read,
                                                   Medipix_sopc_burst_5_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_5_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_5_upstream_write,
                                                   Medipix_sopc_burst_5_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream,
                                                   d1_Medipix_sopc_burst_5_upstream_end_xfer
                                                )
;

  output  [ 26: 0] Medipix_sopc_burst_5_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_5_upstream_burstcount;
  output  [ 28: 0] Medipix_sopc_burst_5_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_5_upstream_byteenable;
  output           Medipix_sopc_burst_5_upstream_debugaccess;
  output           Medipix_sopc_burst_5_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_5_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_5_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_5_upstream_write;
  output  [ 31: 0] Medipix_sopc_burst_5_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream;
  output           d1_Medipix_sopc_burst_5_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_5_upstream_readdata;
  input            Medipix_sopc_burst_5_upstream_readdatavalid;
  input            Medipix_sopc_burst_5_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [ 26: 0] Medipix_sopc_burst_5_upstream_address;
  wire             Medipix_sopc_burst_5_upstream_allgrants;
  wire             Medipix_sopc_burst_5_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_5_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_5_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_5_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_5_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_5_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_5_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_5_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_burstcount;
  wire             Medipix_sopc_burst_5_upstream_burstcount_fifo_empty;
  wire    [ 28: 0] Medipix_sopc_burst_5_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_5_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_5_upstream_debugaccess;
  wire             Medipix_sopc_burst_5_upstream_end_xfer;
  wire             Medipix_sopc_burst_5_upstream_firsttransfer;
  wire             Medipix_sopc_burst_5_upstream_grant_vector;
  wire             Medipix_sopc_burst_5_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_5_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_5_upstream_load_fifo;
  wire             Medipix_sopc_burst_5_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_5_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_5_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_next_burst_count;
  wire             Medipix_sopc_burst_5_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_5_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_5_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_5_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_5_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_5_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_5_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_5_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_5_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_5_upstream_waits_for_read;
  wire             Medipix_sopc_burst_5_upstream_waits_for_write;
  wire             Medipix_sopc_burst_5_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_5_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_5_upstream;
  reg              d1_Medipix_sopc_burst_5_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_5_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_5_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_5_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_5_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream));
  //assign Medipix_sopc_burst_5_upstream_readdatavalid_from_sa = Medipix_sopc_burst_5_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_readdatavalid_from_sa = Medipix_sopc_burst_5_upstream_readdatavalid;

  //assign Medipix_sopc_burst_5_upstream_readdata_from_sa = Medipix_sopc_burst_5_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_readdata_from_sa = Medipix_sopc_burst_5_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream = ({cpu_linux_data_master_address_to_slave[27] , 27'b0} == 28'h0) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_5_upstream_waitrequest_from_sa = Medipix_sopc_burst_5_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_waitrequest_from_sa = Medipix_sopc_burst_5_upstream_waitrequest;

  //Medipix_sopc_burst_5_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_5_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_5_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_5_upstream;

  //Medipix_sopc_burst_5_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_arb_share_counter_next_value = Medipix_sopc_burst_5_upstream_firsttransfer ? (Medipix_sopc_burst_5_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_5_upstream_arb_share_counter ? (Medipix_sopc_burst_5_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_5_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_allgrants = |Medipix_sopc_burst_5_upstream_grant_vector;

  //Medipix_sopc_burst_5_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_end_xfer = ~(Medipix_sopc_burst_5_upstream_waits_for_read | Medipix_sopc_burst_5_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream = Medipix_sopc_burst_5_upstream_end_xfer & (~Medipix_sopc_burst_5_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_5_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream & Medipix_sopc_burst_5_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream & ~Medipix_sopc_burst_5_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_5_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_5_upstream_arb_counter_enable)
          Medipix_sopc_burst_5_upstream_arb_share_counter <= Medipix_sopc_burst_5_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_5_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_5_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_5_upstream & ~Medipix_sopc_burst_5_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_5_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_5_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_5/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_5_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_5_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_5_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_5/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_5_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_5_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_5_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_move_on_to_next_transaction = Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_5_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_5_upstream, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_5_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_5_upstream_module burstcount_fifo_for_Medipix_sopc_burst_5_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_5_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_5_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_5_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read & Medipix_sopc_burst_5_upstream_load_fifo & ~(Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_5_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_5_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_current_burst_minus_one = Medipix_sopc_burst_5_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_5_upstream, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read) & ~Medipix_sopc_burst_5_upstream_load_fifo))? Medipix_sopc_burst_5_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read & Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_5_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_5_upstream_selected_burstcount :
    (Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_5_upstream_transaction_burst_count :
    Medipix_sopc_burst_5_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_5_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_5_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_5_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read)))
          Medipix_sopc_burst_5_upstream_current_burst <= Medipix_sopc_burst_5_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_5_upstream_load_fifo = (~Medipix_sopc_burst_5_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read) & Medipix_sopc_burst_5_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_5_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read) & ~Medipix_sopc_burst_5_upstream_load_fifo | Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_5_upstream_load_fifo <= p0_Medipix_sopc_burst_5_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_5_upstream, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_5_upstream_current_burst_minus_one) & Medipix_sopc_burst_5_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_5_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_5_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_5_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_5_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_5_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_5_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_5_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_5_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream = Medipix_sopc_burst_5_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_5_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_5/upstream, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_5/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_5_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream;

  //allow new arb cycle for Medipix_sopc_burst_5/upstream, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_5_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_5_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_5_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_firsttransfer = Medipix_sopc_burst_5_upstream_begins_xfer ? Medipix_sopc_burst_5_upstream_unreg_firsttransfer : Medipix_sopc_burst_5_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_5_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_5_upstream_slavearbiterlockenable & Medipix_sopc_burst_5_upstream_any_continuerequest);

  //Medipix_sopc_burst_5_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_5_upstream_begins_xfer)
          Medipix_sopc_burst_5_upstream_reg_firsttransfer <= Medipix_sopc_burst_5_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_5_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_5_upstream_write) && (Medipix_sopc_burst_5_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_5_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_5_upstream_read) && (Medipix_sopc_burst_5_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_5_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_5_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_5_upstream_begins_xfer)
          Medipix_sopc_burst_5_upstream_bbt_burstcounter <= Medipix_sopc_burst_5_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_5_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_beginbursttransfer_internal = Medipix_sopc_burst_5_upstream_begins_xfer & (Medipix_sopc_burst_5_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_5_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_5_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream & cpu_linux_data_master_write;

  //Medipix_sopc_burst_5_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_address = cpu_linux_data_master_address_to_slave;

  //d1_Medipix_sopc_burst_5_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_5_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_5_upstream_end_xfer <= Medipix_sopc_burst_5_upstream_end_xfer;
    end


  //Medipix_sopc_burst_5_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_waits_for_read = Medipix_sopc_burst_5_upstream_in_a_read_cycle & Medipix_sopc_burst_5_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_5_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_5_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_5_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_waits_for_write = Medipix_sopc_burst_5_upstream_in_a_write_cycle & Medipix_sopc_burst_5_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_5_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_5_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_5_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_5_upstream_counter = 0;
  //Medipix_sopc_burst_5_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_5_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_5/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_5/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_5_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_5_downstream_address,
                                                     Medipix_sopc_burst_5_downstream_burstcount,
                                                     Medipix_sopc_burst_5_downstream_byteenable,
                                                     Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1,
                                                     Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1,
                                                     Medipix_sopc_burst_5_downstream_read,
                                                     Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1,
                                                     Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register,
                                                     Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1,
                                                     Medipix_sopc_burst_5_downstream_write,
                                                     Medipix_sopc_burst_5_downstream_writedata,
                                                     clk,
                                                     clock_crossing_s1_readdata_from_sa,
                                                     clock_crossing_s1_waitrequest_from_sa,
                                                     d1_clock_crossing_s1_end_xfer,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_5_downstream_address_to_slave,
                                                     Medipix_sopc_burst_5_downstream_latency_counter,
                                                     Medipix_sopc_burst_5_downstream_readdata,
                                                     Medipix_sopc_burst_5_downstream_readdatavalid,
                                                     Medipix_sopc_burst_5_downstream_reset_n,
                                                     Medipix_sopc_burst_5_downstream_waitrequest
                                                  )
;

  output  [ 26: 0] Medipix_sopc_burst_5_downstream_address_to_slave;
  output           Medipix_sopc_burst_5_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_5_downstream_readdata;
  output           Medipix_sopc_burst_5_downstream_readdatavalid;
  output           Medipix_sopc_burst_5_downstream_reset_n;
  output           Medipix_sopc_burst_5_downstream_waitrequest;
  input   [ 26: 0] Medipix_sopc_burst_5_downstream_address;
  input            Medipix_sopc_burst_5_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_5_downstream_byteenable;
  input            Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1;
  input            Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1;
  input            Medipix_sopc_burst_5_downstream_read;
  input            Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1;
  input            Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register;
  input            Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1;
  input            Medipix_sopc_burst_5_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_5_downstream_writedata;
  input            clk;
  input   [ 31: 0] clock_crossing_s1_readdata_from_sa;
  input            clock_crossing_s1_waitrequest_from_sa;
  input            d1_clock_crossing_s1_end_xfer;
  input            reset_n;

  reg     [ 26: 0] Medipix_sopc_burst_5_downstream_address_last_time;
  wire    [ 26: 0] Medipix_sopc_burst_5_downstream_address_to_slave;
  reg              Medipix_sopc_burst_5_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_5_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_5_downstream_is_granted_some_slave;
  reg              Medipix_sopc_burst_5_downstream_latency_counter;
  reg              Medipix_sopc_burst_5_downstream_read_but_no_slave_selected;
  reg              Medipix_sopc_burst_5_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_5_downstream_readdata;
  wire             Medipix_sopc_burst_5_downstream_readdatavalid;
  wire             Medipix_sopc_burst_5_downstream_reset_n;
  wire             Medipix_sopc_burst_5_downstream_run;
  wire             Medipix_sopc_burst_5_downstream_waitrequest;
  reg              Medipix_sopc_burst_5_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_5_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_Medipix_sopc_burst_5_downstream_latency_counter;
  wire             pre_flush_Medipix_sopc_burst_5_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1 | ~Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1) & (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 | ~Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1) & ((~Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1 | ~(Medipix_sopc_burst_5_downstream_read | Medipix_sopc_burst_5_downstream_write) | (1 & ~clock_crossing_s1_waitrequest_from_sa & (Medipix_sopc_burst_5_downstream_read | Medipix_sopc_burst_5_downstream_write)))) & ((~Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1 | ~(Medipix_sopc_burst_5_downstream_read | Medipix_sopc_burst_5_downstream_write) | (1 & ~clock_crossing_s1_waitrequest_from_sa & (Medipix_sopc_burst_5_downstream_read | Medipix_sopc_burst_5_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_5_downstream_address_to_slave = Medipix_sopc_burst_5_downstream_address;

  //Medipix_sopc_burst_5_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_read_but_no_slave_selected <= 0;
      else 
        Medipix_sopc_burst_5_downstream_read_but_no_slave_selected <= Medipix_sopc_burst_5_downstream_read & Medipix_sopc_burst_5_downstream_run & ~Medipix_sopc_burst_5_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign Medipix_sopc_burst_5_downstream_is_granted_some_slave = Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_5_downstream_readdatavalid = Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_5_downstream_readdatavalid = Medipix_sopc_burst_5_downstream_read_but_no_slave_selected |
    pre_flush_Medipix_sopc_burst_5_downstream_readdatavalid;

  //Medipix_sopc_burst_5/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_5_downstream_readdata = clock_crossing_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_waitrequest = ~Medipix_sopc_burst_5_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_latency_counter <= 0;
      else 
        Medipix_sopc_burst_5_downstream_latency_counter <= p1_Medipix_sopc_burst_5_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_Medipix_sopc_burst_5_downstream_latency_counter = ((Medipix_sopc_burst_5_downstream_run & Medipix_sopc_burst_5_downstream_read))? latency_load_value :
    (Medipix_sopc_burst_5_downstream_latency_counter)? Medipix_sopc_burst_5_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //Medipix_sopc_burst_5_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_5_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_5_downstream_address_last_time <= Medipix_sopc_burst_5_downstream_address;
    end


  //Medipix_sopc_burst_5/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_5_downstream_waitrequest & (Medipix_sopc_burst_5_downstream_read | Medipix_sopc_burst_5_downstream_write);
    end


  //Medipix_sopc_burst_5_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_5_downstream_address != Medipix_sopc_burst_5_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_5_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_5_downstream_burstcount_last_time <= Medipix_sopc_burst_5_downstream_burstcount;
    end


  //Medipix_sopc_burst_5_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_5_downstream_burstcount != Medipix_sopc_burst_5_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_5_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_5_downstream_byteenable_last_time <= Medipix_sopc_burst_5_downstream_byteenable;
    end


  //Medipix_sopc_burst_5_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_5_downstream_byteenable != Medipix_sopc_burst_5_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_5_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_5_downstream_read_last_time <= Medipix_sopc_burst_5_downstream_read;
    end


  //Medipix_sopc_burst_5_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_5_downstream_read != Medipix_sopc_burst_5_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_5_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_5_downstream_write_last_time <= Medipix_sopc_burst_5_downstream_write;
    end


  //Medipix_sopc_burst_5_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_5_downstream_write != Medipix_sopc_burst_5_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_5_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_5_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_5_downstream_writedata_last_time <= Medipix_sopc_burst_5_downstream_writedata;
    end


  //Medipix_sopc_burst_5_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_5_downstream_writedata != Medipix_sopc_burst_5_downstream_writedata_last_time) & Medipix_sopc_burst_5_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_5_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_6_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_6_upstream_module (
                                                                                           // inputs:
                                                                                            clear_fifo,
                                                                                            clk,
                                                                                            data_in,
                                                                                            read,
                                                                                            reset_n,
                                                                                            sync_reset,
                                                                                            write,

                                                                                           // outputs:
                                                                                            data_out,
                                                                                            empty,
                                                                                            fifo_contains_ones_n,
                                                                                            full
                                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_6_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_6_upstream_readdata,
                                                   Medipix_sopc_burst_6_upstream_readdatavalid,
                                                   Medipix_sopc_burst_6_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_instruction_master_address_to_slave,
                                                   cpu_linux_instruction_master_burstcount,
                                                   cpu_linux_instruction_master_latency_counter,
                                                   cpu_linux_instruction_master_read,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_6_upstream_address,
                                                   Medipix_sopc_burst_6_upstream_byteaddress,
                                                   Medipix_sopc_burst_6_upstream_byteenable,
                                                   Medipix_sopc_burst_6_upstream_debugaccess,
                                                   Medipix_sopc_burst_6_upstream_read,
                                                   Medipix_sopc_burst_6_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_6_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_6_upstream_write,
                                                   cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream,
                                                   cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream,
                                                   cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register,
                                                   cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream,
                                                   d1_Medipix_sopc_burst_6_upstream_end_xfer
                                                )
;

  output  [ 10: 0] Medipix_sopc_burst_6_upstream_address;
  output  [ 12: 0] Medipix_sopc_burst_6_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_6_upstream_byteenable;
  output           Medipix_sopc_burst_6_upstream_debugaccess;
  output           Medipix_sopc_burst_6_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_6_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_6_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_6_upstream_write;
  output           cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream;
  output           cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream;
  output           cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream;
  output           cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register;
  output           cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream;
  output           d1_Medipix_sopc_burst_6_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_6_upstream_readdata;
  input            Medipix_sopc_burst_6_upstream_readdatavalid;
  input            Medipix_sopc_burst_6_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_instruction_master_address_to_slave;
  input   [  3: 0] cpu_linux_instruction_master_burstcount;
  input            cpu_linux_instruction_master_latency_counter;
  input            cpu_linux_instruction_master_read;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register;
  input            reset_n;

  wire    [ 10: 0] Medipix_sopc_burst_6_upstream_address;
  wire             Medipix_sopc_burst_6_upstream_allgrants;
  wire             Medipix_sopc_burst_6_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_6_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_6_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_6_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_6_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_arb_share_set_values;
  wire             Medipix_sopc_burst_6_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_6_upstream_begins_xfer;
  wire             Medipix_sopc_burst_6_upstream_burstcount_fifo_empty;
  wire    [ 12: 0] Medipix_sopc_burst_6_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_6_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_6_upstream_debugaccess;
  wire             Medipix_sopc_burst_6_upstream_end_xfer;
  wire             Medipix_sopc_burst_6_upstream_firsttransfer;
  wire             Medipix_sopc_burst_6_upstream_grant_vector;
  wire             Medipix_sopc_burst_6_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_6_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_6_upstream_load_fifo;
  wire             Medipix_sopc_burst_6_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_6_upstream_move_on_to_next_transaction;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_next_burst_count;
  wire             Medipix_sopc_burst_6_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_6_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_6_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_6_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_6_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_6_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_6_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_6_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_6_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_6_upstream_waits_for_read;
  wire             Medipix_sopc_burst_6_upstream_waits_for_write;
  wire             Medipix_sopc_burst_6_upstream_write;
  wire             cpu_linux_instruction_master_arbiterlock;
  wire             cpu_linux_instruction_master_arbiterlock2;
  wire             cpu_linux_instruction_master_continuerequest;
  wire             cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_rdv_fifo_output_from_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register;
  wire             cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_6_upstream;
  reg              d1_Medipix_sopc_burst_6_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_6_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_6_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_6_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_6_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream));
  //assign Medipix_sopc_burst_6_upstream_readdatavalid_from_sa = Medipix_sopc_burst_6_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_readdatavalid_from_sa = Medipix_sopc_burst_6_upstream_readdatavalid;

  //assign Medipix_sopc_burst_6_upstream_readdata_from_sa = Medipix_sopc_burst_6_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_readdata_from_sa = Medipix_sopc_burst_6_upstream_readdata;

  assign cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream = (({cpu_linux_instruction_master_address_to_slave[27 : 11] , 11'b0} == 28'h8001800) & (cpu_linux_instruction_master_read)) & cpu_linux_instruction_master_read;
  //assign Medipix_sopc_burst_6_upstream_waitrequest_from_sa = Medipix_sopc_burst_6_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_waitrequest_from_sa = Medipix_sopc_burst_6_upstream_waitrequest;

  //Medipix_sopc_burst_6_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_arb_share_set_values = 1;

  //Medipix_sopc_burst_6_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_6_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_any_bursting_master_saved_grant = cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_6_upstream;

  //Medipix_sopc_burst_6_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_arb_share_counter_next_value = Medipix_sopc_burst_6_upstream_firsttransfer ? (Medipix_sopc_burst_6_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_6_upstream_arb_share_counter ? (Medipix_sopc_burst_6_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_6_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_allgrants = |Medipix_sopc_burst_6_upstream_grant_vector;

  //Medipix_sopc_burst_6_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_end_xfer = ~(Medipix_sopc_burst_6_upstream_waits_for_read | Medipix_sopc_burst_6_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream = Medipix_sopc_burst_6_upstream_end_xfer & (~Medipix_sopc_burst_6_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_6_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream & Medipix_sopc_burst_6_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream & ~Medipix_sopc_burst_6_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_6_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_6_upstream_arb_counter_enable)
          Medipix_sopc_burst_6_upstream_arb_share_counter <= Medipix_sopc_burst_6_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_6_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_6_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_6_upstream & ~Medipix_sopc_burst_6_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_6_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_6_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/instruction_master Medipix_sopc_burst_6/upstream arbiterlock, which is an e_assign
  assign cpu_linux_instruction_master_arbiterlock = Medipix_sopc_burst_6_upstream_slavearbiterlockenable & cpu_linux_instruction_master_continuerequest;

  //Medipix_sopc_burst_6_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_6_upstream_arb_share_counter_next_value;

  //cpu_linux/instruction_master Medipix_sopc_burst_6/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_instruction_master_arbiterlock2 = Medipix_sopc_burst_6_upstream_slavearbiterlockenable2 & cpu_linux_instruction_master_continuerequest;

  //Medipix_sopc_burst_6_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_any_continuerequest = 1;

  //cpu_linux_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_instruction_master_continuerequest = 1;

  assign cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream = cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream & ~((cpu_linux_instruction_master_read & ((cpu_linux_instruction_master_latency_counter != 0) | (1 < cpu_linux_instruction_master_latency_counter) | (|cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register) | (|cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_6_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_move_on_to_next_transaction = Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_6_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_6_upstream, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_selected_burstcount = (cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream)? cpu_linux_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_6_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_6_upstream_module burstcount_fifo_for_Medipix_sopc_burst_6_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_6_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_6_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_6_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read & Medipix_sopc_burst_6_upstream_load_fifo & ~(Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_6_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_6_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_current_burst_minus_one = Medipix_sopc_burst_6_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_6_upstream, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read) & ~Medipix_sopc_burst_6_upstream_load_fifo))? Medipix_sopc_burst_6_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read & Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_6_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_6_upstream_selected_burstcount :
    (Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_6_upstream_transaction_burst_count :
    Medipix_sopc_burst_6_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_6_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_6_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_6_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read)))
          Medipix_sopc_burst_6_upstream_current_burst <= Medipix_sopc_burst_6_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_6_upstream_load_fifo = (~Medipix_sopc_burst_6_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read) & Medipix_sopc_burst_6_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_6_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read) & ~Medipix_sopc_burst_6_upstream_load_fifo | Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_6_upstream_load_fifo <= p0_Medipix_sopc_burst_6_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_6_upstream, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_6_upstream_current_burst_minus_one) & Medipix_sopc_burst_6_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_6_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_6_upstream_module rdv_fifo_for_cpu_linux_instruction_master_to_Medipix_sopc_burst_6_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream),
      .data_out             (cpu_linux_instruction_master_rdv_fifo_output_from_Medipix_sopc_burst_6_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_6_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_6_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_6_upstream_waits_for_read)
    );

  assign cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register = ~cpu_linux_instruction_master_rdv_fifo_empty_Medipix_sopc_burst_6_upstream;
  //local readdatavalid cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream, which is an e_mux
  assign cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream = Medipix_sopc_burst_6_upstream_readdatavalid_from_sa;

  //byteaddress mux for Medipix_sopc_burst_6/upstream, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_byteaddress = cpu_linux_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream = cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream;

  //cpu_linux/instruction_master saved-grant Medipix_sopc_burst_6/upstream, which is an e_assign
  assign cpu_linux_instruction_master_saved_grant_Medipix_sopc_burst_6_upstream = cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream;

  //allow new arb cycle for Medipix_sopc_burst_6/upstream, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_6_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_6_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_6_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_firsttransfer = Medipix_sopc_burst_6_upstream_begins_xfer ? Medipix_sopc_burst_6_upstream_unreg_firsttransfer : Medipix_sopc_burst_6_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_6_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_6_upstream_slavearbiterlockenable & Medipix_sopc_burst_6_upstream_any_continuerequest);

  //Medipix_sopc_burst_6_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_6_upstream_begins_xfer)
          Medipix_sopc_burst_6_upstream_reg_firsttransfer <= Medipix_sopc_burst_6_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_6_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_beginbursttransfer_internal = Medipix_sopc_burst_6_upstream_begins_xfer;

  //Medipix_sopc_burst_6_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_read = cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream & cpu_linux_instruction_master_read;

  //Medipix_sopc_burst_6_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_write = 0;

  //Medipix_sopc_burst_6_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_address = cpu_linux_instruction_master_address_to_slave;

  //d1_Medipix_sopc_burst_6_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_6_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_6_upstream_end_xfer <= Medipix_sopc_burst_6_upstream_end_xfer;
    end


  //Medipix_sopc_burst_6_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_waits_for_read = Medipix_sopc_burst_6_upstream_in_a_read_cycle & Medipix_sopc_burst_6_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_6_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_in_a_read_cycle = cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream & cpu_linux_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_6_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_6_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_waits_for_write = Medipix_sopc_burst_6_upstream_in_a_write_cycle & Medipix_sopc_burst_6_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_6_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_6_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_6_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_6_upstream_counter = 0;
  //Medipix_sopc_burst_6_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_6_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_6/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream && (cpu_linux_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/instruction_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_6/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_6_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_6_downstream_address,
                                                     Medipix_sopc_burst_6_downstream_burstcount,
                                                     Medipix_sopc_burst_6_downstream_byteenable,
                                                     Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_6_downstream_read,
                                                     Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_6_downstream_write,
                                                     Medipix_sopc_burst_6_downstream_writedata,
                                                     clk,
                                                     d1_epcs_controller_epcs_control_port_end_xfer,
                                                     epcs_controller_epcs_control_port_readdata_from_sa,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_6_downstream_address_to_slave,
                                                     Medipix_sopc_burst_6_downstream_latency_counter,
                                                     Medipix_sopc_burst_6_downstream_readdata,
                                                     Medipix_sopc_burst_6_downstream_readdatavalid,
                                                     Medipix_sopc_burst_6_downstream_reset_n,
                                                     Medipix_sopc_burst_6_downstream_waitrequest
                                                  )
;

  output  [ 10: 0] Medipix_sopc_burst_6_downstream_address_to_slave;
  output           Medipix_sopc_burst_6_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_6_downstream_readdata;
  output           Medipix_sopc_burst_6_downstream_readdatavalid;
  output           Medipix_sopc_burst_6_downstream_reset_n;
  output           Medipix_sopc_burst_6_downstream_waitrequest;
  input   [ 10: 0] Medipix_sopc_burst_6_downstream_address;
  input            Medipix_sopc_burst_6_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_6_downstream_byteenable;
  input            Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_6_downstream_read;
  input            Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_6_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_6_downstream_writedata;
  input            clk;
  input            d1_epcs_controller_epcs_control_port_end_xfer;
  input   [ 31: 0] epcs_controller_epcs_control_port_readdata_from_sa;
  input            reset_n;

  reg     [ 10: 0] Medipix_sopc_burst_6_downstream_address_last_time;
  wire    [ 10: 0] Medipix_sopc_burst_6_downstream_address_to_slave;
  reg              Medipix_sopc_burst_6_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_6_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_6_downstream_is_granted_some_slave;
  reg              Medipix_sopc_burst_6_downstream_latency_counter;
  reg              Medipix_sopc_burst_6_downstream_read_but_no_slave_selected;
  reg              Medipix_sopc_burst_6_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_6_downstream_readdata;
  wire             Medipix_sopc_burst_6_downstream_readdatavalid;
  wire             Medipix_sopc_burst_6_downstream_reset_n;
  wire             Medipix_sopc_burst_6_downstream_run;
  wire             Medipix_sopc_burst_6_downstream_waitrequest;
  reg              Medipix_sopc_burst_6_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_6_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_Medipix_sopc_burst_6_downstream_latency_counter;
  wire             pre_flush_Medipix_sopc_burst_6_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port | ~Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port) & (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port | ~Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port) & ((~Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port | ~(Medipix_sopc_burst_6_downstream_read | Medipix_sopc_burst_6_downstream_write) | (1 & ~d1_epcs_controller_epcs_control_port_end_xfer & (Medipix_sopc_burst_6_downstream_read | Medipix_sopc_burst_6_downstream_write)))) & ((~Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port | ~(Medipix_sopc_burst_6_downstream_read | Medipix_sopc_burst_6_downstream_write) | (1 & ~d1_epcs_controller_epcs_control_port_end_xfer & (Medipix_sopc_burst_6_downstream_read | Medipix_sopc_burst_6_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_6_downstream_address_to_slave = Medipix_sopc_burst_6_downstream_address;

  //Medipix_sopc_burst_6_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_read_but_no_slave_selected <= 0;
      else 
        Medipix_sopc_burst_6_downstream_read_but_no_slave_selected <= Medipix_sopc_burst_6_downstream_read & Medipix_sopc_burst_6_downstream_run & ~Medipix_sopc_burst_6_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign Medipix_sopc_burst_6_downstream_is_granted_some_slave = Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_6_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_6_downstream_readdatavalid = Medipix_sopc_burst_6_downstream_read_but_no_slave_selected |
    pre_flush_Medipix_sopc_burst_6_downstream_readdatavalid |
    Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port;

  //Medipix_sopc_burst_6/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_6_downstream_readdata = epcs_controller_epcs_control_port_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_waitrequest = ~Medipix_sopc_burst_6_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_latency_counter <= 0;
      else 
        Medipix_sopc_burst_6_downstream_latency_counter <= p1_Medipix_sopc_burst_6_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_Medipix_sopc_burst_6_downstream_latency_counter = ((Medipix_sopc_burst_6_downstream_run & Medipix_sopc_burst_6_downstream_read))? latency_load_value :
    (Medipix_sopc_burst_6_downstream_latency_counter)? Medipix_sopc_burst_6_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //Medipix_sopc_burst_6_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_6_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_6_downstream_address_last_time <= Medipix_sopc_burst_6_downstream_address;
    end


  //Medipix_sopc_burst_6/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_6_downstream_waitrequest & (Medipix_sopc_burst_6_downstream_read | Medipix_sopc_burst_6_downstream_write);
    end


  //Medipix_sopc_burst_6_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_6_downstream_address != Medipix_sopc_burst_6_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_6_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_6_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_6_downstream_burstcount_last_time <= Medipix_sopc_burst_6_downstream_burstcount;
    end


  //Medipix_sopc_burst_6_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_6_downstream_burstcount != Medipix_sopc_burst_6_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_6_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_6_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_6_downstream_byteenable_last_time <= Medipix_sopc_burst_6_downstream_byteenable;
    end


  //Medipix_sopc_burst_6_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_6_downstream_byteenable != Medipix_sopc_burst_6_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_6_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_6_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_6_downstream_read_last_time <= Medipix_sopc_burst_6_downstream_read;
    end


  //Medipix_sopc_burst_6_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_6_downstream_read != Medipix_sopc_burst_6_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_6_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_6_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_6_downstream_write_last_time <= Medipix_sopc_burst_6_downstream_write;
    end


  //Medipix_sopc_burst_6_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_6_downstream_write != Medipix_sopc_burst_6_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_6_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_6_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_6_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_6_downstream_writedata_last_time <= Medipix_sopc_burst_6_downstream_writedata;
    end


  //Medipix_sopc_burst_6_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_6_downstream_writedata != Medipix_sopc_burst_6_downstream_writedata_last_time) & Medipix_sopc_burst_6_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_6_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_7_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_7_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_7_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_7_upstream_readdata,
                                                   Medipix_sopc_burst_7_upstream_readdatavalid,
                                                   Medipix_sopc_burst_7_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_7_upstream_address,
                                                   Medipix_sopc_burst_7_upstream_burstcount,
                                                   Medipix_sopc_burst_7_upstream_byteaddress,
                                                   Medipix_sopc_burst_7_upstream_byteenable,
                                                   Medipix_sopc_burst_7_upstream_debugaccess,
                                                   Medipix_sopc_burst_7_upstream_read,
                                                   Medipix_sopc_burst_7_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_7_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_7_upstream_write,
                                                   Medipix_sopc_burst_7_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream,
                                                   d1_Medipix_sopc_burst_7_upstream_end_xfer
                                                )
;

  output  [ 10: 0] Medipix_sopc_burst_7_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_7_upstream_burstcount;
  output  [ 12: 0] Medipix_sopc_burst_7_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_7_upstream_byteenable;
  output           Medipix_sopc_burst_7_upstream_debugaccess;
  output           Medipix_sopc_burst_7_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_7_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_7_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_7_upstream_write;
  output  [ 31: 0] Medipix_sopc_burst_7_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream;
  output           d1_Medipix_sopc_burst_7_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_7_upstream_readdata;
  input            Medipix_sopc_burst_7_upstream_readdatavalid;
  input            Medipix_sopc_burst_7_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [ 10: 0] Medipix_sopc_burst_7_upstream_address;
  wire             Medipix_sopc_burst_7_upstream_allgrants;
  wire             Medipix_sopc_burst_7_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_7_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_7_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_7_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_7_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_7_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_7_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_7_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_burstcount;
  wire             Medipix_sopc_burst_7_upstream_burstcount_fifo_empty;
  wire    [ 12: 0] Medipix_sopc_burst_7_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_7_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_7_upstream_debugaccess;
  wire             Medipix_sopc_burst_7_upstream_end_xfer;
  wire             Medipix_sopc_burst_7_upstream_firsttransfer;
  wire             Medipix_sopc_burst_7_upstream_grant_vector;
  wire             Medipix_sopc_burst_7_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_7_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_7_upstream_load_fifo;
  wire             Medipix_sopc_burst_7_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_7_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_7_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_next_burst_count;
  wire             Medipix_sopc_burst_7_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_7_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_7_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_7_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_7_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_7_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_7_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_7_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_7_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_7_upstream_waits_for_read;
  wire             Medipix_sopc_burst_7_upstream_waits_for_write;
  wire             Medipix_sopc_burst_7_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_7_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_7_upstream;
  reg              d1_Medipix_sopc_burst_7_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_7_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_7_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_7_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_7_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream));
  //assign Medipix_sopc_burst_7_upstream_readdatavalid_from_sa = Medipix_sopc_burst_7_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_readdatavalid_from_sa = Medipix_sopc_burst_7_upstream_readdatavalid;

  //assign Medipix_sopc_burst_7_upstream_readdata_from_sa = Medipix_sopc_burst_7_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_readdata_from_sa = Medipix_sopc_burst_7_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream = ({cpu_linux_data_master_address_to_slave[27 : 11] , 11'b0} == 28'h8001800) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_7_upstream_waitrequest_from_sa = Medipix_sopc_burst_7_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_waitrequest_from_sa = Medipix_sopc_burst_7_upstream_waitrequest;

  //Medipix_sopc_burst_7_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_7_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_7_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_7_upstream;

  //Medipix_sopc_burst_7_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_arb_share_counter_next_value = Medipix_sopc_burst_7_upstream_firsttransfer ? (Medipix_sopc_burst_7_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_7_upstream_arb_share_counter ? (Medipix_sopc_burst_7_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_7_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_allgrants = |Medipix_sopc_burst_7_upstream_grant_vector;

  //Medipix_sopc_burst_7_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_end_xfer = ~(Medipix_sopc_burst_7_upstream_waits_for_read | Medipix_sopc_burst_7_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream = Medipix_sopc_burst_7_upstream_end_xfer & (~Medipix_sopc_burst_7_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_7_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream & Medipix_sopc_burst_7_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream & ~Medipix_sopc_burst_7_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_7_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_7_upstream_arb_counter_enable)
          Medipix_sopc_burst_7_upstream_arb_share_counter <= Medipix_sopc_burst_7_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_7_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_7_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_7_upstream & ~Medipix_sopc_burst_7_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_7_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_7_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_7/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_7_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_7_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_7_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_7/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_7_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_7_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_7_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_move_on_to_next_transaction = Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_7_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_7_upstream, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_7_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_7_upstream_module burstcount_fifo_for_Medipix_sopc_burst_7_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_7_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_7_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_7_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read & Medipix_sopc_burst_7_upstream_load_fifo & ~(Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_7_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_7_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_current_burst_minus_one = Medipix_sopc_burst_7_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_7_upstream, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read) & ~Medipix_sopc_burst_7_upstream_load_fifo))? Medipix_sopc_burst_7_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read & Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_7_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_7_upstream_selected_burstcount :
    (Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_7_upstream_transaction_burst_count :
    Medipix_sopc_burst_7_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_7_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_7_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_7_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read)))
          Medipix_sopc_burst_7_upstream_current_burst <= Medipix_sopc_burst_7_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_7_upstream_load_fifo = (~Medipix_sopc_burst_7_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read) & Medipix_sopc_burst_7_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_7_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read) & ~Medipix_sopc_burst_7_upstream_load_fifo | Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_7_upstream_load_fifo <= p0_Medipix_sopc_burst_7_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_7_upstream, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_7_upstream_current_burst_minus_one) & Medipix_sopc_burst_7_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_7_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_7_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_7_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_7_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_7_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_7_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_7_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_7_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream = Medipix_sopc_burst_7_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_7_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_7/upstream, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_7/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_7_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream;

  //allow new arb cycle for Medipix_sopc_burst_7/upstream, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_7_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_7_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_7_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_firsttransfer = Medipix_sopc_burst_7_upstream_begins_xfer ? Medipix_sopc_burst_7_upstream_unreg_firsttransfer : Medipix_sopc_burst_7_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_7_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_7_upstream_slavearbiterlockenable & Medipix_sopc_burst_7_upstream_any_continuerequest);

  //Medipix_sopc_burst_7_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_7_upstream_begins_xfer)
          Medipix_sopc_burst_7_upstream_reg_firsttransfer <= Medipix_sopc_burst_7_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_7_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_7_upstream_write) && (Medipix_sopc_burst_7_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_7_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_7_upstream_read) && (Medipix_sopc_burst_7_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_7_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_7_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_7_upstream_begins_xfer)
          Medipix_sopc_burst_7_upstream_bbt_burstcounter <= Medipix_sopc_burst_7_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_7_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_beginbursttransfer_internal = Medipix_sopc_burst_7_upstream_begins_xfer & (Medipix_sopc_burst_7_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_7_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_7_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream & cpu_linux_data_master_write;

  //Medipix_sopc_burst_7_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_address = cpu_linux_data_master_address_to_slave;

  //d1_Medipix_sopc_burst_7_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_7_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_7_upstream_end_xfer <= Medipix_sopc_burst_7_upstream_end_xfer;
    end


  //Medipix_sopc_burst_7_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_waits_for_read = Medipix_sopc_burst_7_upstream_in_a_read_cycle & Medipix_sopc_burst_7_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_7_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_7_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_7_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_waits_for_write = Medipix_sopc_burst_7_upstream_in_a_write_cycle & Medipix_sopc_burst_7_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_7_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_7_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_7_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_7_upstream_counter = 0;
  //Medipix_sopc_burst_7_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_7_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_7/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_7/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_7_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_7_downstream_address,
                                                     Medipix_sopc_burst_7_downstream_burstcount,
                                                     Medipix_sopc_burst_7_downstream_byteenable,
                                                     Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_7_downstream_read,
                                                     Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port,
                                                     Medipix_sopc_burst_7_downstream_write,
                                                     Medipix_sopc_burst_7_downstream_writedata,
                                                     clk,
                                                     d1_epcs_controller_epcs_control_port_end_xfer,
                                                     epcs_controller_epcs_control_port_readdata_from_sa,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_7_downstream_address_to_slave,
                                                     Medipix_sopc_burst_7_downstream_latency_counter,
                                                     Medipix_sopc_burst_7_downstream_readdata,
                                                     Medipix_sopc_burst_7_downstream_readdatavalid,
                                                     Medipix_sopc_burst_7_downstream_reset_n,
                                                     Medipix_sopc_burst_7_downstream_waitrequest
                                                  )
;

  output  [ 10: 0] Medipix_sopc_burst_7_downstream_address_to_slave;
  output           Medipix_sopc_burst_7_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_7_downstream_readdata;
  output           Medipix_sopc_burst_7_downstream_readdatavalid;
  output           Medipix_sopc_burst_7_downstream_reset_n;
  output           Medipix_sopc_burst_7_downstream_waitrequest;
  input   [ 10: 0] Medipix_sopc_burst_7_downstream_address;
  input            Medipix_sopc_burst_7_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_7_downstream_byteenable;
  input            Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_7_downstream_read;
  input            Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port;
  input            Medipix_sopc_burst_7_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_7_downstream_writedata;
  input            clk;
  input            d1_epcs_controller_epcs_control_port_end_xfer;
  input   [ 31: 0] epcs_controller_epcs_control_port_readdata_from_sa;
  input            reset_n;

  reg     [ 10: 0] Medipix_sopc_burst_7_downstream_address_last_time;
  wire    [ 10: 0] Medipix_sopc_burst_7_downstream_address_to_slave;
  reg              Medipix_sopc_burst_7_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_7_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_7_downstream_is_granted_some_slave;
  reg              Medipix_sopc_burst_7_downstream_latency_counter;
  reg              Medipix_sopc_burst_7_downstream_read_but_no_slave_selected;
  reg              Medipix_sopc_burst_7_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_7_downstream_readdata;
  wire             Medipix_sopc_burst_7_downstream_readdatavalid;
  wire             Medipix_sopc_burst_7_downstream_reset_n;
  wire             Medipix_sopc_burst_7_downstream_run;
  wire             Medipix_sopc_burst_7_downstream_waitrequest;
  reg              Medipix_sopc_burst_7_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_7_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_Medipix_sopc_burst_7_downstream_latency_counter;
  wire             pre_flush_Medipix_sopc_burst_7_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port | ~Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port) & (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port | ~Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port) & ((~Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port | ~(Medipix_sopc_burst_7_downstream_read | Medipix_sopc_burst_7_downstream_write) | (1 & ~d1_epcs_controller_epcs_control_port_end_xfer & (Medipix_sopc_burst_7_downstream_read | Medipix_sopc_burst_7_downstream_write)))) & ((~Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port | ~(Medipix_sopc_burst_7_downstream_read | Medipix_sopc_burst_7_downstream_write) | (1 & ~d1_epcs_controller_epcs_control_port_end_xfer & (Medipix_sopc_burst_7_downstream_read | Medipix_sopc_burst_7_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_7_downstream_address_to_slave = Medipix_sopc_burst_7_downstream_address;

  //Medipix_sopc_burst_7_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_read_but_no_slave_selected <= 0;
      else 
        Medipix_sopc_burst_7_downstream_read_but_no_slave_selected <= Medipix_sopc_burst_7_downstream_read & Medipix_sopc_burst_7_downstream_run & ~Medipix_sopc_burst_7_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign Medipix_sopc_burst_7_downstream_is_granted_some_slave = Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_7_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_7_downstream_readdatavalid = Medipix_sopc_burst_7_downstream_read_but_no_slave_selected |
    pre_flush_Medipix_sopc_burst_7_downstream_readdatavalid |
    Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port;

  //Medipix_sopc_burst_7/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_7_downstream_readdata = epcs_controller_epcs_control_port_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_waitrequest = ~Medipix_sopc_burst_7_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_latency_counter <= 0;
      else 
        Medipix_sopc_burst_7_downstream_latency_counter <= p1_Medipix_sopc_burst_7_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_Medipix_sopc_burst_7_downstream_latency_counter = ((Medipix_sopc_burst_7_downstream_run & Medipix_sopc_burst_7_downstream_read))? latency_load_value :
    (Medipix_sopc_burst_7_downstream_latency_counter)? Medipix_sopc_burst_7_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //Medipix_sopc_burst_7_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_7_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_7_downstream_address_last_time <= Medipix_sopc_burst_7_downstream_address;
    end


  //Medipix_sopc_burst_7/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_7_downstream_waitrequest & (Medipix_sopc_burst_7_downstream_read | Medipix_sopc_burst_7_downstream_write);
    end


  //Medipix_sopc_burst_7_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_7_downstream_address != Medipix_sopc_burst_7_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_7_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_7_downstream_burstcount_last_time <= Medipix_sopc_burst_7_downstream_burstcount;
    end


  //Medipix_sopc_burst_7_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_7_downstream_burstcount != Medipix_sopc_burst_7_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_7_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_7_downstream_byteenable_last_time <= Medipix_sopc_burst_7_downstream_byteenable;
    end


  //Medipix_sopc_burst_7_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_7_downstream_byteenable != Medipix_sopc_burst_7_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_7_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_7_downstream_read_last_time <= Medipix_sopc_burst_7_downstream_read;
    end


  //Medipix_sopc_burst_7_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_7_downstream_read != Medipix_sopc_burst_7_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_7_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_7_downstream_write_last_time <= Medipix_sopc_burst_7_downstream_write;
    end


  //Medipix_sopc_burst_7_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_7_downstream_write != Medipix_sopc_burst_7_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_7_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_7_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_7_downstream_writedata_last_time <= Medipix_sopc_burst_7_downstream_writedata;
    end


  //Medipix_sopc_burst_7_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_7_downstream_writedata != Medipix_sopc_burst_7_downstream_writedata_last_time) & Medipix_sopc_burst_7_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_7_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_8_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_8_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_8_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_8_upstream_readdata,
                                                   Medipix_sopc_burst_8_upstream_readdatavalid,
                                                   Medipix_sopc_burst_8_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_8_upstream_address,
                                                   Medipix_sopc_burst_8_upstream_burstcount,
                                                   Medipix_sopc_burst_8_upstream_byteaddress,
                                                   Medipix_sopc_burst_8_upstream_byteenable,
                                                   Medipix_sopc_burst_8_upstream_debugaccess,
                                                   Medipix_sopc_burst_8_upstream_read,
                                                   Medipix_sopc_burst_8_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_8_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_8_upstream_write,
                                                   Medipix_sopc_burst_8_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream,
                                                   d1_Medipix_sopc_burst_8_upstream_end_xfer
                                                )
;

  output  [ 11: 0] Medipix_sopc_burst_8_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_8_upstream_burstcount;
  output  [ 13: 0] Medipix_sopc_burst_8_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_8_upstream_byteenable;
  output           Medipix_sopc_burst_8_upstream_debugaccess;
  output           Medipix_sopc_burst_8_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_8_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_8_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_8_upstream_write;
  output  [ 31: 0] Medipix_sopc_burst_8_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream;
  output           d1_Medipix_sopc_burst_8_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_8_upstream_readdata;
  input            Medipix_sopc_burst_8_upstream_readdatavalid;
  input            Medipix_sopc_burst_8_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [ 11: 0] Medipix_sopc_burst_8_upstream_address;
  wire             Medipix_sopc_burst_8_upstream_allgrants;
  wire             Medipix_sopc_burst_8_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_8_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_8_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_8_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_8_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_8_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_8_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_8_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_burstcount;
  wire             Medipix_sopc_burst_8_upstream_burstcount_fifo_empty;
  wire    [ 13: 0] Medipix_sopc_burst_8_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_8_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_8_upstream_debugaccess;
  wire             Medipix_sopc_burst_8_upstream_end_xfer;
  wire             Medipix_sopc_burst_8_upstream_firsttransfer;
  wire             Medipix_sopc_burst_8_upstream_grant_vector;
  wire             Medipix_sopc_burst_8_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_8_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_8_upstream_load_fifo;
  wire             Medipix_sopc_burst_8_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_8_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_8_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_next_burst_count;
  wire             Medipix_sopc_burst_8_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_8_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_8_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_8_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_8_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_8_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_8_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_8_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_8_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_8_upstream_waits_for_read;
  wire             Medipix_sopc_burst_8_upstream_waits_for_write;
  wire             Medipix_sopc_burst_8_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_8_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_8_upstream;
  reg              d1_Medipix_sopc_burst_8_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_8_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_8_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_8_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_8_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream));
  //assign Medipix_sopc_burst_8_upstream_readdatavalid_from_sa = Medipix_sopc_burst_8_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_readdatavalid_from_sa = Medipix_sopc_burst_8_upstream_readdatavalid;

  //assign Medipix_sopc_burst_8_upstream_readdata_from_sa = Medipix_sopc_burst_8_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_readdata_from_sa = Medipix_sopc_burst_8_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream = ({cpu_linux_data_master_address_to_slave[27 : 12] , 12'b0} == 28'h8002000) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_8_upstream_waitrequest_from_sa = Medipix_sopc_burst_8_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_waitrequest_from_sa = Medipix_sopc_burst_8_upstream_waitrequest;

  //Medipix_sopc_burst_8_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_8_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_8_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_8_upstream;

  //Medipix_sopc_burst_8_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_arb_share_counter_next_value = Medipix_sopc_burst_8_upstream_firsttransfer ? (Medipix_sopc_burst_8_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_8_upstream_arb_share_counter ? (Medipix_sopc_burst_8_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_8_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_allgrants = |Medipix_sopc_burst_8_upstream_grant_vector;

  //Medipix_sopc_burst_8_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_end_xfer = ~(Medipix_sopc_burst_8_upstream_waits_for_read | Medipix_sopc_burst_8_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream = Medipix_sopc_burst_8_upstream_end_xfer & (~Medipix_sopc_burst_8_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_8_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream & Medipix_sopc_burst_8_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream & ~Medipix_sopc_burst_8_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_8_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_8_upstream_arb_counter_enable)
          Medipix_sopc_burst_8_upstream_arb_share_counter <= Medipix_sopc_burst_8_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_8_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_8_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_8_upstream & ~Medipix_sopc_burst_8_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_8_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_8_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_8/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_8_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_8_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_8_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_8/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_8_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_8_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_8_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_move_on_to_next_transaction = Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_8_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_8_upstream, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_8_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_8_upstream_module burstcount_fifo_for_Medipix_sopc_burst_8_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_8_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_8_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_8_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read & Medipix_sopc_burst_8_upstream_load_fifo & ~(Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_8_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_8_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_current_burst_minus_one = Medipix_sopc_burst_8_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_8_upstream, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read) & ~Medipix_sopc_burst_8_upstream_load_fifo))? Medipix_sopc_burst_8_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read & Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_8_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_8_upstream_selected_burstcount :
    (Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_8_upstream_transaction_burst_count :
    Medipix_sopc_burst_8_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_8_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_8_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_8_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read)))
          Medipix_sopc_burst_8_upstream_current_burst <= Medipix_sopc_burst_8_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_8_upstream_load_fifo = (~Medipix_sopc_burst_8_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read) & Medipix_sopc_burst_8_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_8_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read) & ~Medipix_sopc_burst_8_upstream_load_fifo | Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_8_upstream_load_fifo <= p0_Medipix_sopc_burst_8_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_8_upstream, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_8_upstream_current_burst_minus_one) & Medipix_sopc_burst_8_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_8_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_8_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_8_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_8_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_8_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_8_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_8_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_8_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream = Medipix_sopc_burst_8_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_8_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_8/upstream, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_8/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_8_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream;

  //allow new arb cycle for Medipix_sopc_burst_8/upstream, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_8_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_8_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_8_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_firsttransfer = Medipix_sopc_burst_8_upstream_begins_xfer ? Medipix_sopc_burst_8_upstream_unreg_firsttransfer : Medipix_sopc_burst_8_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_8_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_8_upstream_slavearbiterlockenable & Medipix_sopc_burst_8_upstream_any_continuerequest);

  //Medipix_sopc_burst_8_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_8_upstream_begins_xfer)
          Medipix_sopc_burst_8_upstream_reg_firsttransfer <= Medipix_sopc_burst_8_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_8_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_8_upstream_write) && (Medipix_sopc_burst_8_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_8_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_8_upstream_read) && (Medipix_sopc_burst_8_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_8_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_8_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_8_upstream_begins_xfer)
          Medipix_sopc_burst_8_upstream_bbt_burstcounter <= Medipix_sopc_burst_8_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_8_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_beginbursttransfer_internal = Medipix_sopc_burst_8_upstream_begins_xfer & (Medipix_sopc_burst_8_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_8_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_8_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream & cpu_linux_data_master_write;

  //Medipix_sopc_burst_8_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_address = cpu_linux_data_master_address_to_slave;

  //d1_Medipix_sopc_burst_8_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_8_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_8_upstream_end_xfer <= Medipix_sopc_burst_8_upstream_end_xfer;
    end


  //Medipix_sopc_burst_8_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_waits_for_read = Medipix_sopc_burst_8_upstream_in_a_read_cycle & Medipix_sopc_burst_8_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_8_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_8_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_8_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_waits_for_write = Medipix_sopc_burst_8_upstream_in_a_write_cycle & Medipix_sopc_burst_8_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_8_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_8_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_8_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_8_upstream_counter = 0;
  //Medipix_sopc_burst_8_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_8_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_8/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_8/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_8_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_8_downstream_address,
                                                     Medipix_sopc_burst_8_downstream_burstcount,
                                                     Medipix_sopc_burst_8_downstream_byteenable,
                                                     Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port,
                                                     Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port,
                                                     Medipix_sopc_burst_8_downstream_read,
                                                     Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port,
                                                     Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port,
                                                     Medipix_sopc_burst_8_downstream_write,
                                                     Medipix_sopc_burst_8_downstream_writedata,
                                                     clk,
                                                     d1_igor_mac_control_port_end_xfer,
                                                     igor_mac_control_port_readdata_from_sa,
                                                     igor_mac_control_port_waitrequest_n_from_sa,
                                                     reset_n,

                                                    // outputs:
                                                     Medipix_sopc_burst_8_downstream_address_to_slave,
                                                     Medipix_sopc_burst_8_downstream_latency_counter,
                                                     Medipix_sopc_burst_8_downstream_readdata,
                                                     Medipix_sopc_burst_8_downstream_readdatavalid,
                                                     Medipix_sopc_burst_8_downstream_reset_n,
                                                     Medipix_sopc_burst_8_downstream_waitrequest
                                                  )
;

  output  [ 11: 0] Medipix_sopc_burst_8_downstream_address_to_slave;
  output           Medipix_sopc_burst_8_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_8_downstream_readdata;
  output           Medipix_sopc_burst_8_downstream_readdatavalid;
  output           Medipix_sopc_burst_8_downstream_reset_n;
  output           Medipix_sopc_burst_8_downstream_waitrequest;
  input   [ 11: 0] Medipix_sopc_burst_8_downstream_address;
  input            Medipix_sopc_burst_8_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_8_downstream_byteenable;
  input            Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port;
  input            Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port;
  input            Medipix_sopc_burst_8_downstream_read;
  input            Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port;
  input            Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port;
  input            Medipix_sopc_burst_8_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_8_downstream_writedata;
  input            clk;
  input            d1_igor_mac_control_port_end_xfer;
  input   [ 31: 0] igor_mac_control_port_readdata_from_sa;
  input            igor_mac_control_port_waitrequest_n_from_sa;
  input            reset_n;

  reg     [ 11: 0] Medipix_sopc_burst_8_downstream_address_last_time;
  wire    [ 11: 0] Medipix_sopc_burst_8_downstream_address_to_slave;
  reg              Medipix_sopc_burst_8_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_8_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_8_downstream_latency_counter;
  reg              Medipix_sopc_burst_8_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_8_downstream_readdata;
  wire             Medipix_sopc_burst_8_downstream_readdatavalid;
  wire             Medipix_sopc_burst_8_downstream_reset_n;
  wire             Medipix_sopc_burst_8_downstream_run;
  wire             Medipix_sopc_burst_8_downstream_waitrequest;
  reg              Medipix_sopc_burst_8_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_8_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             pre_flush_Medipix_sopc_burst_8_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port | ~Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port) & ((~Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port | ~(Medipix_sopc_burst_8_downstream_read | Medipix_sopc_burst_8_downstream_write) | (1 & igor_mac_control_port_waitrequest_n_from_sa & (Medipix_sopc_burst_8_downstream_read | Medipix_sopc_burst_8_downstream_write)))) & ((~Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port | ~(Medipix_sopc_burst_8_downstream_read | Medipix_sopc_burst_8_downstream_write) | (1 & igor_mac_control_port_waitrequest_n_from_sa & (Medipix_sopc_burst_8_downstream_read | Medipix_sopc_burst_8_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_8_downstream_address_to_slave = Medipix_sopc_burst_8_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_8_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_8_downstream_readdatavalid = 0 |
    pre_flush_Medipix_sopc_burst_8_downstream_readdatavalid |
    Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port;

  //Medipix_sopc_burst_8/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_8_downstream_readdata = igor_mac_control_port_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_waitrequest = ~Medipix_sopc_burst_8_downstream_run;

  //latent max counter, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_latency_counter = 0;

  //Medipix_sopc_burst_8_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_8_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_8_downstream_address_last_time <= Medipix_sopc_burst_8_downstream_address;
    end


  //Medipix_sopc_burst_8/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_8_downstream_waitrequest & (Medipix_sopc_burst_8_downstream_read | Medipix_sopc_burst_8_downstream_write);
    end


  //Medipix_sopc_burst_8_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_8_downstream_address != Medipix_sopc_burst_8_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_8_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_8_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_8_downstream_burstcount_last_time <= Medipix_sopc_burst_8_downstream_burstcount;
    end


  //Medipix_sopc_burst_8_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_8_downstream_burstcount != Medipix_sopc_burst_8_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_8_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_8_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_8_downstream_byteenable_last_time <= Medipix_sopc_burst_8_downstream_byteenable;
    end


  //Medipix_sopc_burst_8_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_8_downstream_byteenable != Medipix_sopc_burst_8_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_8_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_8_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_8_downstream_read_last_time <= Medipix_sopc_burst_8_downstream_read;
    end


  //Medipix_sopc_burst_8_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_8_downstream_read != Medipix_sopc_burst_8_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_8_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_8_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_8_downstream_write_last_time <= Medipix_sopc_burst_8_downstream_write;
    end


  //Medipix_sopc_burst_8_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_8_downstream_write != Medipix_sopc_burst_8_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_8_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_8_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_8_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_8_downstream_writedata_last_time <= Medipix_sopc_burst_8_downstream_writedata;
    end


  //Medipix_sopc_burst_8_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_8_downstream_writedata != Medipix_sopc_burst_8_downstream_writedata_last_time) & Medipix_sopc_burst_8_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_8_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_Medipix_sopc_burst_9_upstream_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_9_upstream_module (
                                                                                    // inputs:
                                                                                     clear_fifo,
                                                                                     clk,
                                                                                     data_in,
                                                                                     read,
                                                                                     reset_n,
                                                                                     sync_reset,
                                                                                     write,

                                                                                    // outputs:
                                                                                     data_out,
                                                                                     empty,
                                                                                     fifo_contains_ones_n,
                                                                                     full
                                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_9_upstream_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_9_upstream_readdata,
                                                   Medipix_sopc_burst_9_upstream_readdatavalid,
                                                   Medipix_sopc_burst_9_upstream_waitrequest,
                                                   clk,
                                                   cpu_linux_data_master_address_to_slave,
                                                   cpu_linux_data_master_burstcount,
                                                   cpu_linux_data_master_byteenable,
                                                   cpu_linux_data_master_debugaccess,
                                                   cpu_linux_data_master_latency_counter,
                                                   cpu_linux_data_master_read,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                                   cpu_linux_data_master_write,
                                                   cpu_linux_data_master_writedata,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_9_upstream_address,
                                                   Medipix_sopc_burst_9_upstream_burstcount,
                                                   Medipix_sopc_burst_9_upstream_byteaddress,
                                                   Medipix_sopc_burst_9_upstream_byteenable,
                                                   Medipix_sopc_burst_9_upstream_debugaccess,
                                                   Medipix_sopc_burst_9_upstream_read,
                                                   Medipix_sopc_burst_9_upstream_readdata_from_sa,
                                                   Medipix_sopc_burst_9_upstream_waitrequest_from_sa,
                                                   Medipix_sopc_burst_9_upstream_write,
                                                   Medipix_sopc_burst_9_upstream_writedata,
                                                   cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream,
                                                   cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream,
                                                   cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                                   cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream,
                                                   d1_Medipix_sopc_burst_9_upstream_end_xfer
                                                )
;

  output  [  3: 0] Medipix_sopc_burst_9_upstream_address;
  output  [  3: 0] Medipix_sopc_burst_9_upstream_burstcount;
  output  [  5: 0] Medipix_sopc_burst_9_upstream_byteaddress;
  output  [  3: 0] Medipix_sopc_burst_9_upstream_byteenable;
  output           Medipix_sopc_burst_9_upstream_debugaccess;
  output           Medipix_sopc_burst_9_upstream_read;
  output  [ 31: 0] Medipix_sopc_burst_9_upstream_readdata_from_sa;
  output           Medipix_sopc_burst_9_upstream_waitrequest_from_sa;
  output           Medipix_sopc_burst_9_upstream_write;
  output  [ 31: 0] Medipix_sopc_burst_9_upstream_writedata;
  output           cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream;
  output           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream;
  output           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  output           cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream;
  output           d1_Medipix_sopc_burst_9_upstream_end_xfer;
  input   [ 31: 0] Medipix_sopc_burst_9_upstream_readdata;
  input            Medipix_sopc_burst_9_upstream_readdatavalid;
  input            Medipix_sopc_burst_9_upstream_waitrequest;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address_to_slave;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_debugaccess;
  input            cpu_linux_data_master_latency_counter;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            reset_n;

  wire    [  3: 0] Medipix_sopc_burst_9_upstream_address;
  wire             Medipix_sopc_burst_9_upstream_allgrants;
  wire             Medipix_sopc_burst_9_upstream_allow_new_arb_cycle;
  wire             Medipix_sopc_burst_9_upstream_any_bursting_master_saved_grant;
  wire             Medipix_sopc_burst_9_upstream_any_continuerequest;
  wire             Medipix_sopc_burst_9_upstream_arb_counter_enable;
  reg     [  3: 0] Medipix_sopc_burst_9_upstream_arb_share_counter;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_arb_share_counter_next_value;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_arb_share_set_values;
  reg     [  2: 0] Medipix_sopc_burst_9_upstream_bbt_burstcounter;
  wire             Medipix_sopc_burst_9_upstream_beginbursttransfer_internal;
  wire             Medipix_sopc_burst_9_upstream_begins_xfer;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_burstcount;
  wire             Medipix_sopc_burst_9_upstream_burstcount_fifo_empty;
  wire    [  5: 0] Medipix_sopc_burst_9_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_byteenable;
  reg     [  3: 0] Medipix_sopc_burst_9_upstream_current_burst;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_current_burst_minus_one;
  wire             Medipix_sopc_burst_9_upstream_debugaccess;
  wire             Medipix_sopc_burst_9_upstream_end_xfer;
  wire             Medipix_sopc_burst_9_upstream_firsttransfer;
  wire             Medipix_sopc_burst_9_upstream_grant_vector;
  wire             Medipix_sopc_burst_9_upstream_in_a_read_cycle;
  wire             Medipix_sopc_burst_9_upstream_in_a_write_cycle;
  reg              Medipix_sopc_burst_9_upstream_load_fifo;
  wire             Medipix_sopc_burst_9_upstream_master_qreq_vector;
  wire             Medipix_sopc_burst_9_upstream_move_on_to_next_transaction;
  wire    [  2: 0] Medipix_sopc_burst_9_upstream_next_bbt_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_next_burst_count;
  wire             Medipix_sopc_burst_9_upstream_non_bursting_master_requests;
  wire             Medipix_sopc_burst_9_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_9_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_9_upstream_readdatavalid_from_sa;
  reg              Medipix_sopc_burst_9_upstream_reg_firsttransfer;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_selected_burstcount;
  reg              Medipix_sopc_burst_9_upstream_slavearbiterlockenable;
  wire             Medipix_sopc_burst_9_upstream_slavearbiterlockenable2;
  wire             Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_transaction_burst_count;
  wire             Medipix_sopc_burst_9_upstream_unreg_firsttransfer;
  wire             Medipix_sopc_burst_9_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_9_upstream_waits_for_read;
  wire             Medipix_sopc_burst_9_upstream_waits_for_write;
  wire             Medipix_sopc_burst_9_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_9_upstream_writedata;
  wire             cpu_linux_data_master_arbiterlock;
  wire             cpu_linux_data_master_arbiterlock2;
  wire             cpu_linux_data_master_continuerequest;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_saved_grant_Medipix_sopc_burst_9_upstream;
  reg              d1_Medipix_sopc_burst_9_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_Medipix_sopc_burst_9_upstream_load_fifo;
  wire             wait_for_Medipix_sopc_burst_9_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~Medipix_sopc_burst_9_upstream_end_xfer;
    end


  assign Medipix_sopc_burst_9_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream));
  //assign Medipix_sopc_burst_9_upstream_readdatavalid_from_sa = Medipix_sopc_burst_9_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_readdatavalid_from_sa = Medipix_sopc_burst_9_upstream_readdatavalid;

  //assign Medipix_sopc_burst_9_upstream_readdata_from_sa = Medipix_sopc_burst_9_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_readdata_from_sa = Medipix_sopc_burst_9_upstream_readdata;

  assign cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream = ({cpu_linux_data_master_address_to_slave[27 : 4] , 4'b0} == 28'h8000000) & (cpu_linux_data_master_read | cpu_linux_data_master_write);
  //assign Medipix_sopc_burst_9_upstream_waitrequest_from_sa = Medipix_sopc_burst_9_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_waitrequest_from_sa = Medipix_sopc_burst_9_upstream_waitrequest;

  //Medipix_sopc_burst_9_upstream_arb_share_counter set values, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_arb_share_set_values = (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream)? (((cpu_linux_data_master_write) ? cpu_linux_data_master_burstcount : 1)) :
    1;

  //Medipix_sopc_burst_9_upstream_non_bursting_master_requests mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_non_bursting_master_requests = 0;

  //Medipix_sopc_burst_9_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_any_bursting_master_saved_grant = cpu_linux_data_master_saved_grant_Medipix_sopc_burst_9_upstream;

  //Medipix_sopc_burst_9_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_arb_share_counter_next_value = Medipix_sopc_burst_9_upstream_firsttransfer ? (Medipix_sopc_burst_9_upstream_arb_share_set_values - 1) : |Medipix_sopc_burst_9_upstream_arb_share_counter ? (Medipix_sopc_burst_9_upstream_arb_share_counter - 1) : 0;

  //Medipix_sopc_burst_9_upstream_allgrants all slave grants, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_allgrants = |Medipix_sopc_burst_9_upstream_grant_vector;

  //Medipix_sopc_burst_9_upstream_end_xfer assignment, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_end_xfer = ~(Medipix_sopc_burst_9_upstream_waits_for_read | Medipix_sopc_burst_9_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream = Medipix_sopc_burst_9_upstream_end_xfer & (~Medipix_sopc_burst_9_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //Medipix_sopc_burst_9_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream & Medipix_sopc_burst_9_upstream_allgrants) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream & ~Medipix_sopc_burst_9_upstream_non_bursting_master_requests);

  //Medipix_sopc_burst_9_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_upstream_arb_share_counter <= 0;
      else if (Medipix_sopc_burst_9_upstream_arb_counter_enable)
          Medipix_sopc_burst_9_upstream_arb_share_counter <= Medipix_sopc_burst_9_upstream_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_9_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_upstream_slavearbiterlockenable <= 0;
      else if ((|Medipix_sopc_burst_9_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream) | (end_xfer_arb_share_counter_term_Medipix_sopc_burst_9_upstream & ~Medipix_sopc_burst_9_upstream_non_bursting_master_requests))
          Medipix_sopc_burst_9_upstream_slavearbiterlockenable <= |Medipix_sopc_burst_9_upstream_arb_share_counter_next_value;
    end


  //cpu_linux/data_master Medipix_sopc_burst_9/upstream arbiterlock, which is an e_assign
  assign cpu_linux_data_master_arbiterlock = Medipix_sopc_burst_9_upstream_slavearbiterlockenable & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_9_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_slavearbiterlockenable2 = |Medipix_sopc_burst_9_upstream_arb_share_counter_next_value;

  //cpu_linux/data_master Medipix_sopc_burst_9/upstream arbiterlock2, which is an e_assign
  assign cpu_linux_data_master_arbiterlock2 = Medipix_sopc_burst_9_upstream_slavearbiterlockenable2 & cpu_linux_data_master_continuerequest;

  //Medipix_sopc_burst_9_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_any_continuerequest = 1;

  //cpu_linux_data_master_continuerequest continued request, which is an e_assign
  assign cpu_linux_data_master_continuerequest = 1;

  assign cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream & ~((cpu_linux_data_master_read & ((cpu_linux_data_master_latency_counter != 0) | (1 < cpu_linux_data_master_latency_counter) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register) | (|cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register))));
  //unique name for Medipix_sopc_burst_9_upstream_move_on_to_next_transaction, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_move_on_to_next_transaction = Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_9_upstream_load_fifo;

  //the currently selected burstcount for Medipix_sopc_burst_9_upstream, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_selected_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream)? cpu_linux_data_master_burstcount :
    1;

  //burstcount_fifo_for_Medipix_sopc_burst_9_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_Medipix_sopc_burst_9_upstream_module burstcount_fifo_for_Medipix_sopc_burst_9_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_9_upstream_selected_burstcount),
      .data_out             (Medipix_sopc_burst_9_upstream_transaction_burst_count),
      .empty                (Medipix_sopc_burst_9_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read & Medipix_sopc_burst_9_upstream_load_fifo & ~(Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_9_upstream_burstcount_fifo_empty))
    );

  //Medipix_sopc_burst_9_upstream current burst minus one, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_current_burst_minus_one = Medipix_sopc_burst_9_upstream_current_burst - 1;

  //what to load in current_burst, for Medipix_sopc_burst_9_upstream, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_next_burst_count = (((in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read) & ~Medipix_sopc_burst_9_upstream_load_fifo))? Medipix_sopc_burst_9_upstream_selected_burstcount :
    ((in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read & Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst & Medipix_sopc_burst_9_upstream_burstcount_fifo_empty))? Medipix_sopc_burst_9_upstream_selected_burstcount :
    (Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst)? Medipix_sopc_burst_9_upstream_transaction_burst_count :
    Medipix_sopc_burst_9_upstream_current_burst_minus_one;

  //the current burst count for Medipix_sopc_burst_9_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_upstream_current_burst <= 0;
      else if (Medipix_sopc_burst_9_upstream_readdatavalid_from_sa | (~Medipix_sopc_burst_9_upstream_load_fifo & (in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read)))
          Medipix_sopc_burst_9_upstream_current_burst <= Medipix_sopc_burst_9_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_Medipix_sopc_burst_9_upstream_load_fifo = (~Medipix_sopc_burst_9_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read) & Medipix_sopc_burst_9_upstream_load_fifo))? 1 :
    ~Medipix_sopc_burst_9_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read) & ~Medipix_sopc_burst_9_upstream_load_fifo | Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst)
          Medipix_sopc_burst_9_upstream_load_fifo <= p0_Medipix_sopc_burst_9_upstream_load_fifo;
    end


  //the last cycle in the burst for Medipix_sopc_burst_9_upstream, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_this_cycle_is_the_last_burst = ~(|Medipix_sopc_burst_9_upstream_current_burst_minus_one) & Medipix_sopc_burst_9_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_9_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_9_upstream_module rdv_fifo_for_cpu_linux_data_master_to_Medipix_sopc_burst_9_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream),
      .data_out             (cpu_linux_data_master_rdv_fifo_output_from_Medipix_sopc_burst_9_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_9_upstream),
      .full                 (),
      .read                 (Medipix_sopc_burst_9_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~Medipix_sopc_burst_9_upstream_waits_for_read)
    );

  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register = ~cpu_linux_data_master_rdv_fifo_empty_Medipix_sopc_burst_9_upstream;
  //local readdatavalid cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream, which is an e_mux
  assign cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream = Medipix_sopc_burst_9_upstream_readdatavalid_from_sa;

  //Medipix_sopc_burst_9_upstream_writedata mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_writedata = cpu_linux_data_master_writedata;

  //byteaddress mux for Medipix_sopc_burst_9/upstream, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_byteaddress = cpu_linux_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream = cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream;

  //cpu_linux/data_master saved-grant Medipix_sopc_burst_9/upstream, which is an e_assign
  assign cpu_linux_data_master_saved_grant_Medipix_sopc_burst_9_upstream = cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream;

  //allow new arb cycle for Medipix_sopc_burst_9/upstream, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign Medipix_sopc_burst_9_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign Medipix_sopc_burst_9_upstream_master_qreq_vector = 1;

  //Medipix_sopc_burst_9_upstream_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_firsttransfer = Medipix_sopc_burst_9_upstream_begins_xfer ? Medipix_sopc_burst_9_upstream_unreg_firsttransfer : Medipix_sopc_burst_9_upstream_reg_firsttransfer;

  //Medipix_sopc_burst_9_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_unreg_firsttransfer = ~(Medipix_sopc_burst_9_upstream_slavearbiterlockenable & Medipix_sopc_burst_9_upstream_any_continuerequest);

  //Medipix_sopc_burst_9_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_upstream_reg_firsttransfer <= 1'b1;
      else if (Medipix_sopc_burst_9_upstream_begins_xfer)
          Medipix_sopc_burst_9_upstream_reg_firsttransfer <= Medipix_sopc_burst_9_upstream_unreg_firsttransfer;
    end


  //Medipix_sopc_burst_9_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_next_bbt_burstcount = ((((Medipix_sopc_burst_9_upstream_write) && (Medipix_sopc_burst_9_upstream_bbt_burstcounter == 0))))? (Medipix_sopc_burst_9_upstream_burstcount - 1) :
    ((((Medipix_sopc_burst_9_upstream_read) && (Medipix_sopc_burst_9_upstream_bbt_burstcounter == 0))))? 0 :
    (Medipix_sopc_burst_9_upstream_bbt_burstcounter - 1);

  //Medipix_sopc_burst_9_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_upstream_bbt_burstcounter <= 0;
      else if (Medipix_sopc_burst_9_upstream_begins_xfer)
          Medipix_sopc_burst_9_upstream_bbt_burstcounter <= Medipix_sopc_burst_9_upstream_next_bbt_burstcount;
    end


  //Medipix_sopc_burst_9_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_beginbursttransfer_internal = Medipix_sopc_burst_9_upstream_begins_xfer & (Medipix_sopc_burst_9_upstream_bbt_burstcounter == 0);

  //Medipix_sopc_burst_9_upstream_read assignment, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_read = cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream & cpu_linux_data_master_read;

  //Medipix_sopc_burst_9_upstream_write assignment, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_write = cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream & cpu_linux_data_master_write;

  //Medipix_sopc_burst_9_upstream_address mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_address = cpu_linux_data_master_address_to_slave;

  //d1_Medipix_sopc_burst_9_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_Medipix_sopc_burst_9_upstream_end_xfer <= 1;
      else 
        d1_Medipix_sopc_burst_9_upstream_end_xfer <= Medipix_sopc_burst_9_upstream_end_xfer;
    end


  //Medipix_sopc_burst_9_upstream_waits_for_read in a cycle, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_waits_for_read = Medipix_sopc_burst_9_upstream_in_a_read_cycle & Medipix_sopc_burst_9_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_9_upstream_in_a_read_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_in_a_read_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream & cpu_linux_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = Medipix_sopc_burst_9_upstream_in_a_read_cycle;

  //Medipix_sopc_burst_9_upstream_waits_for_write in a cycle, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_waits_for_write = Medipix_sopc_burst_9_upstream_in_a_write_cycle & Medipix_sopc_burst_9_upstream_waitrequest_from_sa;

  //Medipix_sopc_burst_9_upstream_in_a_write_cycle assignment, which is an e_assign
  assign Medipix_sopc_burst_9_upstream_in_a_write_cycle = cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream & cpu_linux_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = Medipix_sopc_burst_9_upstream_in_a_write_cycle;

  assign wait_for_Medipix_sopc_burst_9_upstream_counter = 0;
  //Medipix_sopc_burst_9_upstream_byteenable byte enable port mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_byteenable = (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream)? cpu_linux_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_burstcount = (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream)? cpu_linux_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign Medipix_sopc_burst_9_upstream_debugaccess = (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream)? cpu_linux_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_9/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu_linux/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream && (cpu_linux_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu_linux/data_master drove 0 on its 'burstcount' port while accessing slave Medipix_sopc_burst_9/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_burst_9_downstream_arbitrator (
                                                    // inputs:
                                                     Medipix_sopc_burst_9_downstream_address,
                                                     Medipix_sopc_burst_9_downstream_burstcount,
                                                     Medipix_sopc_burst_9_downstream_byteenable,
                                                     Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0,
                                                     Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0,
                                                     Medipix_sopc_burst_9_downstream_read,
                                                     Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0,
                                                     Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0,
                                                     Medipix_sopc_burst_9_downstream_write,
                                                     Medipix_sopc_burst_9_downstream_writedata,
                                                     clk,
                                                     d1_tx_table_avalon_slave_0_end_xfer,
                                                     reset_n,
                                                     tx_table_avalon_slave_0_readdata_from_sa,

                                                    // outputs:
                                                     Medipix_sopc_burst_9_downstream_address_to_slave,
                                                     Medipix_sopc_burst_9_downstream_latency_counter,
                                                     Medipix_sopc_burst_9_downstream_readdata,
                                                     Medipix_sopc_burst_9_downstream_readdatavalid,
                                                     Medipix_sopc_burst_9_downstream_reset_n,
                                                     Medipix_sopc_burst_9_downstream_waitrequest
                                                  )
;

  output  [  3: 0] Medipix_sopc_burst_9_downstream_address_to_slave;
  output           Medipix_sopc_burst_9_downstream_latency_counter;
  output  [ 31: 0] Medipix_sopc_burst_9_downstream_readdata;
  output           Medipix_sopc_burst_9_downstream_readdatavalid;
  output           Medipix_sopc_burst_9_downstream_reset_n;
  output           Medipix_sopc_burst_9_downstream_waitrequest;
  input   [  3: 0] Medipix_sopc_burst_9_downstream_address;
  input            Medipix_sopc_burst_9_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_9_downstream_byteenable;
  input            Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0;
  input            Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0;
  input            Medipix_sopc_burst_9_downstream_read;
  input            Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0;
  input            Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0;
  input            Medipix_sopc_burst_9_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_9_downstream_writedata;
  input            clk;
  input            d1_tx_table_avalon_slave_0_end_xfer;
  input            reset_n;
  input   [ 31: 0] tx_table_avalon_slave_0_readdata_from_sa;

  reg     [  3: 0] Medipix_sopc_burst_9_downstream_address_last_time;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_address_to_slave;
  reg              Medipix_sopc_burst_9_downstream_burstcount_last_time;
  reg     [  3: 0] Medipix_sopc_burst_9_downstream_byteenable_last_time;
  wire             Medipix_sopc_burst_9_downstream_latency_counter;
  reg              Medipix_sopc_burst_9_downstream_read_last_time;
  wire    [ 31: 0] Medipix_sopc_burst_9_downstream_readdata;
  wire             Medipix_sopc_burst_9_downstream_readdatavalid;
  wire             Medipix_sopc_burst_9_downstream_reset_n;
  wire             Medipix_sopc_burst_9_downstream_run;
  wire             Medipix_sopc_burst_9_downstream_waitrequest;
  reg              Medipix_sopc_burst_9_downstream_write_last_time;
  reg     [ 31: 0] Medipix_sopc_burst_9_downstream_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             pre_flush_Medipix_sopc_burst_9_downstream_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0 | ~Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0) & ((~Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0 | ~Medipix_sopc_burst_9_downstream_read | (1 & ~d1_tx_table_avalon_slave_0_end_xfer & Medipix_sopc_burst_9_downstream_read))) & ((~Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0 | ~Medipix_sopc_burst_9_downstream_write | (1 & Medipix_sopc_burst_9_downstream_write)));

  //cascaded wait assignment, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign Medipix_sopc_burst_9_downstream_address_to_slave = Medipix_sopc_burst_9_downstream_address;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_Medipix_sopc_burst_9_downstream_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign Medipix_sopc_burst_9_downstream_readdatavalid = 0 |
    pre_flush_Medipix_sopc_burst_9_downstream_readdatavalid |
    Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0;

  //Medipix_sopc_burst_9/downstream readdata mux, which is an e_mux
  assign Medipix_sopc_burst_9_downstream_readdata = tx_table_avalon_slave_0_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_waitrequest = ~Medipix_sopc_burst_9_downstream_run;

  //latent max counter, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_latency_counter = 0;

  //Medipix_sopc_burst_9_downstream_reset_n assignment, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Medipix_sopc_burst_9_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_downstream_address_last_time <= 0;
      else 
        Medipix_sopc_burst_9_downstream_address_last_time <= Medipix_sopc_burst_9_downstream_address;
    end


  //Medipix_sopc_burst_9/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= Medipix_sopc_burst_9_downstream_waitrequest & (Medipix_sopc_burst_9_downstream_read | Medipix_sopc_burst_9_downstream_write);
    end


  //Medipix_sopc_burst_9_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_9_downstream_address != Medipix_sopc_burst_9_downstream_address_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_9_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_9_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_downstream_burstcount_last_time <= 0;
      else 
        Medipix_sopc_burst_9_downstream_burstcount_last_time <= Medipix_sopc_burst_9_downstream_burstcount;
    end


  //Medipix_sopc_burst_9_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_9_downstream_burstcount != Medipix_sopc_burst_9_downstream_burstcount_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_9_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_9_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_downstream_byteenable_last_time <= 0;
      else 
        Medipix_sopc_burst_9_downstream_byteenable_last_time <= Medipix_sopc_burst_9_downstream_byteenable;
    end


  //Medipix_sopc_burst_9_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_9_downstream_byteenable != Medipix_sopc_burst_9_downstream_byteenable_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_9_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_9_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_downstream_read_last_time <= 0;
      else 
        Medipix_sopc_burst_9_downstream_read_last_time <= Medipix_sopc_burst_9_downstream_read;
    end


  //Medipix_sopc_burst_9_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_9_downstream_read != Medipix_sopc_burst_9_downstream_read_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_9_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_9_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_downstream_write_last_time <= 0;
      else 
        Medipix_sopc_burst_9_downstream_write_last_time <= Medipix_sopc_burst_9_downstream_write;
    end


  //Medipix_sopc_burst_9_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_9_downstream_write != Medipix_sopc_burst_9_downstream_write_last_time))
        begin
          $write("%0d ns: Medipix_sopc_burst_9_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_9_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          Medipix_sopc_burst_9_downstream_writedata_last_time <= 0;
      else 
        Medipix_sopc_burst_9_downstream_writedata_last_time <= Medipix_sopc_burst_9_downstream_writedata;
    end


  //Medipix_sopc_burst_9_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (Medipix_sopc_burst_9_downstream_writedata != Medipix_sopc_burst_9_downstream_writedata_last_time) & Medipix_sopc_burst_9_downstream_write)
        begin
          $write("%0d ns: Medipix_sopc_burst_9_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_Medipix_sopc_burst_4_downstream_to_clock_crossing_s1_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  wire             full_96;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_95;
  assign empty = !full_0;
  assign full_96 = 0;
  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    0;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_Medipix_sopc_burst_5_downstream_to_clock_crossing_s1_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  wire             full_96;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_95;
  assign empty = !full_0;
  assign full_96 = 0;
  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    0;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_igor_mac_tx_master_to_clock_crossing_s1_module (
                                                                     // inputs:
                                                                      clear_fifo,
                                                                      clk,
                                                                      data_in,
                                                                      read,
                                                                      reset_n,
                                                                      sync_reset,
                                                                      write,

                                                                     // outputs:
                                                                      data_out,
                                                                      empty,
                                                                      fifo_contains_ones_n,
                                                                      full
                                                                   )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  reg              full_54;
  reg              full_55;
  reg              full_56;
  reg              full_57;
  reg              full_58;
  reg              full_59;
  reg              full_6;
  reg              full_60;
  reg              full_61;
  reg              full_62;
  reg              full_63;
  reg              full_64;
  reg              full_65;
  reg              full_66;
  reg              full_67;
  reg              full_68;
  reg              full_69;
  reg              full_7;
  reg              full_70;
  reg              full_71;
  reg              full_72;
  reg              full_73;
  reg              full_74;
  reg              full_75;
  reg              full_76;
  reg              full_77;
  reg              full_78;
  reg              full_79;
  reg              full_8;
  reg              full_80;
  reg              full_81;
  reg              full_82;
  reg              full_83;
  reg              full_84;
  reg              full_85;
  reg              full_86;
  reg              full_87;
  reg              full_88;
  reg              full_89;
  reg              full_9;
  reg              full_90;
  reg              full_91;
  reg              full_92;
  reg              full_93;
  reg              full_94;
  reg              full_95;
  wire             full_96;
  reg     [  7: 0] how_many_ones;
  wire    [  7: 0] one_count_minus_one;
  wire    [  7: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p54_full_54;
  wire             p54_stage_54;
  wire             p55_full_55;
  wire             p55_stage_55;
  wire             p56_full_56;
  wire             p56_stage_56;
  wire             p57_full_57;
  wire             p57_stage_57;
  wire             p58_full_58;
  wire             p58_stage_58;
  wire             p59_full_59;
  wire             p59_stage_59;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p60_full_60;
  wire             p60_stage_60;
  wire             p61_full_61;
  wire             p61_stage_61;
  wire             p62_full_62;
  wire             p62_stage_62;
  wire             p63_full_63;
  wire             p63_stage_63;
  wire             p64_full_64;
  wire             p64_stage_64;
  wire             p65_full_65;
  wire             p65_stage_65;
  wire             p66_full_66;
  wire             p66_stage_66;
  wire             p67_full_67;
  wire             p67_stage_67;
  wire             p68_full_68;
  wire             p68_stage_68;
  wire             p69_full_69;
  wire             p69_stage_69;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p70_full_70;
  wire             p70_stage_70;
  wire             p71_full_71;
  wire             p71_stage_71;
  wire             p72_full_72;
  wire             p72_stage_72;
  wire             p73_full_73;
  wire             p73_stage_73;
  wire             p74_full_74;
  wire             p74_stage_74;
  wire             p75_full_75;
  wire             p75_stage_75;
  wire             p76_full_76;
  wire             p76_stage_76;
  wire             p77_full_77;
  wire             p77_stage_77;
  wire             p78_full_78;
  wire             p78_stage_78;
  wire             p79_full_79;
  wire             p79_stage_79;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p80_full_80;
  wire             p80_stage_80;
  wire             p81_full_81;
  wire             p81_stage_81;
  wire             p82_full_82;
  wire             p82_stage_82;
  wire             p83_full_83;
  wire             p83_stage_83;
  wire             p84_full_84;
  wire             p84_stage_84;
  wire             p85_full_85;
  wire             p85_stage_85;
  wire             p86_full_86;
  wire             p86_stage_86;
  wire             p87_full_87;
  wire             p87_stage_87;
  wire             p88_full_88;
  wire             p88_stage_88;
  wire             p89_full_89;
  wire             p89_stage_89;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p90_full_90;
  wire             p90_stage_90;
  wire             p91_full_91;
  wire             p91_stage_91;
  wire             p92_full_92;
  wire             p92_stage_92;
  wire             p93_full_93;
  wire             p93_stage_93;
  wire             p94_full_94;
  wire             p94_stage_94;
  wire             p95_full_95;
  wire             p95_stage_95;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_54;
  reg              stage_55;
  reg              stage_56;
  reg              stage_57;
  reg              stage_58;
  reg              stage_59;
  reg              stage_6;
  reg              stage_60;
  reg              stage_61;
  reg              stage_62;
  reg              stage_63;
  reg              stage_64;
  reg              stage_65;
  reg              stage_66;
  reg              stage_67;
  reg              stage_68;
  reg              stage_69;
  reg              stage_7;
  reg              stage_70;
  reg              stage_71;
  reg              stage_72;
  reg              stage_73;
  reg              stage_74;
  reg              stage_75;
  reg              stage_76;
  reg              stage_77;
  reg              stage_78;
  reg              stage_79;
  reg              stage_8;
  reg              stage_80;
  reg              stage_81;
  reg              stage_82;
  reg              stage_83;
  reg              stage_84;
  reg              stage_85;
  reg              stage_86;
  reg              stage_87;
  reg              stage_88;
  reg              stage_89;
  reg              stage_9;
  reg              stage_90;
  reg              stage_91;
  reg              stage_92;
  reg              stage_93;
  reg              stage_94;
  reg              stage_95;
  wire    [  7: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_95;
  assign empty = !full_0;
  assign full_96 = 0;
  //data_95, which is an e_mux
  assign p95_stage_95 = ((full_96 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_95 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_95))
          if (sync_reset & full_95 & !((full_96 == 0) & read & write))
              stage_95 <= 0;
          else 
            stage_95 <= p95_stage_95;
    end


  //control_95, which is an e_mux
  assign p95_full_95 = ((read & !write) == 0)? full_94 :
    0;

  //control_reg_95, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_95 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_95 <= 0;
          else 
            full_95 <= p95_full_95;
    end


  //data_94, which is an e_mux
  assign p94_stage_94 = ((full_95 & ~clear_fifo) == 0)? data_in :
    stage_95;

  //data_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_94 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_94))
          if (sync_reset & full_94 & !((full_95 == 0) & read & write))
              stage_94 <= 0;
          else 
            stage_94 <= p94_stage_94;
    end


  //control_94, which is an e_mux
  assign p94_full_94 = ((read & !write) == 0)? full_93 :
    full_95;

  //control_reg_94, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_94 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_94 <= 0;
          else 
            full_94 <= p94_full_94;
    end


  //data_93, which is an e_mux
  assign p93_stage_93 = ((full_94 & ~clear_fifo) == 0)? data_in :
    stage_94;

  //data_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_93 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_93))
          if (sync_reset & full_93 & !((full_94 == 0) & read & write))
              stage_93 <= 0;
          else 
            stage_93 <= p93_stage_93;
    end


  //control_93, which is an e_mux
  assign p93_full_93 = ((read & !write) == 0)? full_92 :
    full_94;

  //control_reg_93, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_93 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_93 <= 0;
          else 
            full_93 <= p93_full_93;
    end


  //data_92, which is an e_mux
  assign p92_stage_92 = ((full_93 & ~clear_fifo) == 0)? data_in :
    stage_93;

  //data_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_92 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_92))
          if (sync_reset & full_92 & !((full_93 == 0) & read & write))
              stage_92 <= 0;
          else 
            stage_92 <= p92_stage_92;
    end


  //control_92, which is an e_mux
  assign p92_full_92 = ((read & !write) == 0)? full_91 :
    full_93;

  //control_reg_92, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_92 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_92 <= 0;
          else 
            full_92 <= p92_full_92;
    end


  //data_91, which is an e_mux
  assign p91_stage_91 = ((full_92 & ~clear_fifo) == 0)? data_in :
    stage_92;

  //data_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_91 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_91))
          if (sync_reset & full_91 & !((full_92 == 0) & read & write))
              stage_91 <= 0;
          else 
            stage_91 <= p91_stage_91;
    end


  //control_91, which is an e_mux
  assign p91_full_91 = ((read & !write) == 0)? full_90 :
    full_92;

  //control_reg_91, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_91 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_91 <= 0;
          else 
            full_91 <= p91_full_91;
    end


  //data_90, which is an e_mux
  assign p90_stage_90 = ((full_91 & ~clear_fifo) == 0)? data_in :
    stage_91;

  //data_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_90 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_90))
          if (sync_reset & full_90 & !((full_91 == 0) & read & write))
              stage_90 <= 0;
          else 
            stage_90 <= p90_stage_90;
    end


  //control_90, which is an e_mux
  assign p90_full_90 = ((read & !write) == 0)? full_89 :
    full_91;

  //control_reg_90, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_90 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_90 <= 0;
          else 
            full_90 <= p90_full_90;
    end


  //data_89, which is an e_mux
  assign p89_stage_89 = ((full_90 & ~clear_fifo) == 0)? data_in :
    stage_90;

  //data_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_89 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_89))
          if (sync_reset & full_89 & !((full_90 == 0) & read & write))
              stage_89 <= 0;
          else 
            stage_89 <= p89_stage_89;
    end


  //control_89, which is an e_mux
  assign p89_full_89 = ((read & !write) == 0)? full_88 :
    full_90;

  //control_reg_89, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_89 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_89 <= 0;
          else 
            full_89 <= p89_full_89;
    end


  //data_88, which is an e_mux
  assign p88_stage_88 = ((full_89 & ~clear_fifo) == 0)? data_in :
    stage_89;

  //data_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_88 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_88))
          if (sync_reset & full_88 & !((full_89 == 0) & read & write))
              stage_88 <= 0;
          else 
            stage_88 <= p88_stage_88;
    end


  //control_88, which is an e_mux
  assign p88_full_88 = ((read & !write) == 0)? full_87 :
    full_89;

  //control_reg_88, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_88 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_88 <= 0;
          else 
            full_88 <= p88_full_88;
    end


  //data_87, which is an e_mux
  assign p87_stage_87 = ((full_88 & ~clear_fifo) == 0)? data_in :
    stage_88;

  //data_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_87 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_87))
          if (sync_reset & full_87 & !((full_88 == 0) & read & write))
              stage_87 <= 0;
          else 
            stage_87 <= p87_stage_87;
    end


  //control_87, which is an e_mux
  assign p87_full_87 = ((read & !write) == 0)? full_86 :
    full_88;

  //control_reg_87, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_87 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_87 <= 0;
          else 
            full_87 <= p87_full_87;
    end


  //data_86, which is an e_mux
  assign p86_stage_86 = ((full_87 & ~clear_fifo) == 0)? data_in :
    stage_87;

  //data_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_86 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_86))
          if (sync_reset & full_86 & !((full_87 == 0) & read & write))
              stage_86 <= 0;
          else 
            stage_86 <= p86_stage_86;
    end


  //control_86, which is an e_mux
  assign p86_full_86 = ((read & !write) == 0)? full_85 :
    full_87;

  //control_reg_86, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_86 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_86 <= 0;
          else 
            full_86 <= p86_full_86;
    end


  //data_85, which is an e_mux
  assign p85_stage_85 = ((full_86 & ~clear_fifo) == 0)? data_in :
    stage_86;

  //data_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_85 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_85))
          if (sync_reset & full_85 & !((full_86 == 0) & read & write))
              stage_85 <= 0;
          else 
            stage_85 <= p85_stage_85;
    end


  //control_85, which is an e_mux
  assign p85_full_85 = ((read & !write) == 0)? full_84 :
    full_86;

  //control_reg_85, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_85 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_85 <= 0;
          else 
            full_85 <= p85_full_85;
    end


  //data_84, which is an e_mux
  assign p84_stage_84 = ((full_85 & ~clear_fifo) == 0)? data_in :
    stage_85;

  //data_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_84 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_84))
          if (sync_reset & full_84 & !((full_85 == 0) & read & write))
              stage_84 <= 0;
          else 
            stage_84 <= p84_stage_84;
    end


  //control_84, which is an e_mux
  assign p84_full_84 = ((read & !write) == 0)? full_83 :
    full_85;

  //control_reg_84, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_84 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_84 <= 0;
          else 
            full_84 <= p84_full_84;
    end


  //data_83, which is an e_mux
  assign p83_stage_83 = ((full_84 & ~clear_fifo) == 0)? data_in :
    stage_84;

  //data_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_83 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_83))
          if (sync_reset & full_83 & !((full_84 == 0) & read & write))
              stage_83 <= 0;
          else 
            stage_83 <= p83_stage_83;
    end


  //control_83, which is an e_mux
  assign p83_full_83 = ((read & !write) == 0)? full_82 :
    full_84;

  //control_reg_83, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_83 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_83 <= 0;
          else 
            full_83 <= p83_full_83;
    end


  //data_82, which is an e_mux
  assign p82_stage_82 = ((full_83 & ~clear_fifo) == 0)? data_in :
    stage_83;

  //data_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_82 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_82))
          if (sync_reset & full_82 & !((full_83 == 0) & read & write))
              stage_82 <= 0;
          else 
            stage_82 <= p82_stage_82;
    end


  //control_82, which is an e_mux
  assign p82_full_82 = ((read & !write) == 0)? full_81 :
    full_83;

  //control_reg_82, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_82 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_82 <= 0;
          else 
            full_82 <= p82_full_82;
    end


  //data_81, which is an e_mux
  assign p81_stage_81 = ((full_82 & ~clear_fifo) == 0)? data_in :
    stage_82;

  //data_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_81 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_81))
          if (sync_reset & full_81 & !((full_82 == 0) & read & write))
              stage_81 <= 0;
          else 
            stage_81 <= p81_stage_81;
    end


  //control_81, which is an e_mux
  assign p81_full_81 = ((read & !write) == 0)? full_80 :
    full_82;

  //control_reg_81, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_81 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_81 <= 0;
          else 
            full_81 <= p81_full_81;
    end


  //data_80, which is an e_mux
  assign p80_stage_80 = ((full_81 & ~clear_fifo) == 0)? data_in :
    stage_81;

  //data_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_80 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_80))
          if (sync_reset & full_80 & !((full_81 == 0) & read & write))
              stage_80 <= 0;
          else 
            stage_80 <= p80_stage_80;
    end


  //control_80, which is an e_mux
  assign p80_full_80 = ((read & !write) == 0)? full_79 :
    full_81;

  //control_reg_80, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_80 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_80 <= 0;
          else 
            full_80 <= p80_full_80;
    end


  //data_79, which is an e_mux
  assign p79_stage_79 = ((full_80 & ~clear_fifo) == 0)? data_in :
    stage_80;

  //data_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_79 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_79))
          if (sync_reset & full_79 & !((full_80 == 0) & read & write))
              stage_79 <= 0;
          else 
            stage_79 <= p79_stage_79;
    end


  //control_79, which is an e_mux
  assign p79_full_79 = ((read & !write) == 0)? full_78 :
    full_80;

  //control_reg_79, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_79 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_79 <= 0;
          else 
            full_79 <= p79_full_79;
    end


  //data_78, which is an e_mux
  assign p78_stage_78 = ((full_79 & ~clear_fifo) == 0)? data_in :
    stage_79;

  //data_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_78 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_78))
          if (sync_reset & full_78 & !((full_79 == 0) & read & write))
              stage_78 <= 0;
          else 
            stage_78 <= p78_stage_78;
    end


  //control_78, which is an e_mux
  assign p78_full_78 = ((read & !write) == 0)? full_77 :
    full_79;

  //control_reg_78, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_78 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_78 <= 0;
          else 
            full_78 <= p78_full_78;
    end


  //data_77, which is an e_mux
  assign p77_stage_77 = ((full_78 & ~clear_fifo) == 0)? data_in :
    stage_78;

  //data_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_77 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_77))
          if (sync_reset & full_77 & !((full_78 == 0) & read & write))
              stage_77 <= 0;
          else 
            stage_77 <= p77_stage_77;
    end


  //control_77, which is an e_mux
  assign p77_full_77 = ((read & !write) == 0)? full_76 :
    full_78;

  //control_reg_77, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_77 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_77 <= 0;
          else 
            full_77 <= p77_full_77;
    end


  //data_76, which is an e_mux
  assign p76_stage_76 = ((full_77 & ~clear_fifo) == 0)? data_in :
    stage_77;

  //data_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_76 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_76))
          if (sync_reset & full_76 & !((full_77 == 0) & read & write))
              stage_76 <= 0;
          else 
            stage_76 <= p76_stage_76;
    end


  //control_76, which is an e_mux
  assign p76_full_76 = ((read & !write) == 0)? full_75 :
    full_77;

  //control_reg_76, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_76 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_76 <= 0;
          else 
            full_76 <= p76_full_76;
    end


  //data_75, which is an e_mux
  assign p75_stage_75 = ((full_76 & ~clear_fifo) == 0)? data_in :
    stage_76;

  //data_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_75 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_75))
          if (sync_reset & full_75 & !((full_76 == 0) & read & write))
              stage_75 <= 0;
          else 
            stage_75 <= p75_stage_75;
    end


  //control_75, which is an e_mux
  assign p75_full_75 = ((read & !write) == 0)? full_74 :
    full_76;

  //control_reg_75, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_75 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_75 <= 0;
          else 
            full_75 <= p75_full_75;
    end


  //data_74, which is an e_mux
  assign p74_stage_74 = ((full_75 & ~clear_fifo) == 0)? data_in :
    stage_75;

  //data_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_74 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_74))
          if (sync_reset & full_74 & !((full_75 == 0) & read & write))
              stage_74 <= 0;
          else 
            stage_74 <= p74_stage_74;
    end


  //control_74, which is an e_mux
  assign p74_full_74 = ((read & !write) == 0)? full_73 :
    full_75;

  //control_reg_74, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_74 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_74 <= 0;
          else 
            full_74 <= p74_full_74;
    end


  //data_73, which is an e_mux
  assign p73_stage_73 = ((full_74 & ~clear_fifo) == 0)? data_in :
    stage_74;

  //data_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_73 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_73))
          if (sync_reset & full_73 & !((full_74 == 0) & read & write))
              stage_73 <= 0;
          else 
            stage_73 <= p73_stage_73;
    end


  //control_73, which is an e_mux
  assign p73_full_73 = ((read & !write) == 0)? full_72 :
    full_74;

  //control_reg_73, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_73 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_73 <= 0;
          else 
            full_73 <= p73_full_73;
    end


  //data_72, which is an e_mux
  assign p72_stage_72 = ((full_73 & ~clear_fifo) == 0)? data_in :
    stage_73;

  //data_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_72 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_72))
          if (sync_reset & full_72 & !((full_73 == 0) & read & write))
              stage_72 <= 0;
          else 
            stage_72 <= p72_stage_72;
    end


  //control_72, which is an e_mux
  assign p72_full_72 = ((read & !write) == 0)? full_71 :
    full_73;

  //control_reg_72, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_72 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_72 <= 0;
          else 
            full_72 <= p72_full_72;
    end


  //data_71, which is an e_mux
  assign p71_stage_71 = ((full_72 & ~clear_fifo) == 0)? data_in :
    stage_72;

  //data_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_71 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_71))
          if (sync_reset & full_71 & !((full_72 == 0) & read & write))
              stage_71 <= 0;
          else 
            stage_71 <= p71_stage_71;
    end


  //control_71, which is an e_mux
  assign p71_full_71 = ((read & !write) == 0)? full_70 :
    full_72;

  //control_reg_71, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_71 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_71 <= 0;
          else 
            full_71 <= p71_full_71;
    end


  //data_70, which is an e_mux
  assign p70_stage_70 = ((full_71 & ~clear_fifo) == 0)? data_in :
    stage_71;

  //data_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_70 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_70))
          if (sync_reset & full_70 & !((full_71 == 0) & read & write))
              stage_70 <= 0;
          else 
            stage_70 <= p70_stage_70;
    end


  //control_70, which is an e_mux
  assign p70_full_70 = ((read & !write) == 0)? full_69 :
    full_71;

  //control_reg_70, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_70 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_70 <= 0;
          else 
            full_70 <= p70_full_70;
    end


  //data_69, which is an e_mux
  assign p69_stage_69 = ((full_70 & ~clear_fifo) == 0)? data_in :
    stage_70;

  //data_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_69 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_69))
          if (sync_reset & full_69 & !((full_70 == 0) & read & write))
              stage_69 <= 0;
          else 
            stage_69 <= p69_stage_69;
    end


  //control_69, which is an e_mux
  assign p69_full_69 = ((read & !write) == 0)? full_68 :
    full_70;

  //control_reg_69, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_69 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_69 <= 0;
          else 
            full_69 <= p69_full_69;
    end


  //data_68, which is an e_mux
  assign p68_stage_68 = ((full_69 & ~clear_fifo) == 0)? data_in :
    stage_69;

  //data_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_68 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_68))
          if (sync_reset & full_68 & !((full_69 == 0) & read & write))
              stage_68 <= 0;
          else 
            stage_68 <= p68_stage_68;
    end


  //control_68, which is an e_mux
  assign p68_full_68 = ((read & !write) == 0)? full_67 :
    full_69;

  //control_reg_68, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_68 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_68 <= 0;
          else 
            full_68 <= p68_full_68;
    end


  //data_67, which is an e_mux
  assign p67_stage_67 = ((full_68 & ~clear_fifo) == 0)? data_in :
    stage_68;

  //data_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_67 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_67))
          if (sync_reset & full_67 & !((full_68 == 0) & read & write))
              stage_67 <= 0;
          else 
            stage_67 <= p67_stage_67;
    end


  //control_67, which is an e_mux
  assign p67_full_67 = ((read & !write) == 0)? full_66 :
    full_68;

  //control_reg_67, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_67 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_67 <= 0;
          else 
            full_67 <= p67_full_67;
    end


  //data_66, which is an e_mux
  assign p66_stage_66 = ((full_67 & ~clear_fifo) == 0)? data_in :
    stage_67;

  //data_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_66 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_66))
          if (sync_reset & full_66 & !((full_67 == 0) & read & write))
              stage_66 <= 0;
          else 
            stage_66 <= p66_stage_66;
    end


  //control_66, which is an e_mux
  assign p66_full_66 = ((read & !write) == 0)? full_65 :
    full_67;

  //control_reg_66, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_66 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_66 <= 0;
          else 
            full_66 <= p66_full_66;
    end


  //data_65, which is an e_mux
  assign p65_stage_65 = ((full_66 & ~clear_fifo) == 0)? data_in :
    stage_66;

  //data_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_65 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_65))
          if (sync_reset & full_65 & !((full_66 == 0) & read & write))
              stage_65 <= 0;
          else 
            stage_65 <= p65_stage_65;
    end


  //control_65, which is an e_mux
  assign p65_full_65 = ((read & !write) == 0)? full_64 :
    full_66;

  //control_reg_65, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_65 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_65 <= 0;
          else 
            full_65 <= p65_full_65;
    end


  //data_64, which is an e_mux
  assign p64_stage_64 = ((full_65 & ~clear_fifo) == 0)? data_in :
    stage_65;

  //data_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_64 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_64))
          if (sync_reset & full_64 & !((full_65 == 0) & read & write))
              stage_64 <= 0;
          else 
            stage_64 <= p64_stage_64;
    end


  //control_64, which is an e_mux
  assign p64_full_64 = ((read & !write) == 0)? full_63 :
    full_65;

  //control_reg_64, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_64 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_64 <= 0;
          else 
            full_64 <= p64_full_64;
    end


  //data_63, which is an e_mux
  assign p63_stage_63 = ((full_64 & ~clear_fifo) == 0)? data_in :
    stage_64;

  //data_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_63 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_63))
          if (sync_reset & full_63 & !((full_64 == 0) & read & write))
              stage_63 <= 0;
          else 
            stage_63 <= p63_stage_63;
    end


  //control_63, which is an e_mux
  assign p63_full_63 = ((read & !write) == 0)? full_62 :
    full_64;

  //control_reg_63, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_63 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_63 <= 0;
          else 
            full_63 <= p63_full_63;
    end


  //data_62, which is an e_mux
  assign p62_stage_62 = ((full_63 & ~clear_fifo) == 0)? data_in :
    stage_63;

  //data_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_62 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_62))
          if (sync_reset & full_62 & !((full_63 == 0) & read & write))
              stage_62 <= 0;
          else 
            stage_62 <= p62_stage_62;
    end


  //control_62, which is an e_mux
  assign p62_full_62 = ((read & !write) == 0)? full_61 :
    full_63;

  //control_reg_62, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_62 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_62 <= 0;
          else 
            full_62 <= p62_full_62;
    end


  //data_61, which is an e_mux
  assign p61_stage_61 = ((full_62 & ~clear_fifo) == 0)? data_in :
    stage_62;

  //data_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_61 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_61))
          if (sync_reset & full_61 & !((full_62 == 0) & read & write))
              stage_61 <= 0;
          else 
            stage_61 <= p61_stage_61;
    end


  //control_61, which is an e_mux
  assign p61_full_61 = ((read & !write) == 0)? full_60 :
    full_62;

  //control_reg_61, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_61 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_61 <= 0;
          else 
            full_61 <= p61_full_61;
    end


  //data_60, which is an e_mux
  assign p60_stage_60 = ((full_61 & ~clear_fifo) == 0)? data_in :
    stage_61;

  //data_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_60 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_60))
          if (sync_reset & full_60 & !((full_61 == 0) & read & write))
              stage_60 <= 0;
          else 
            stage_60 <= p60_stage_60;
    end


  //control_60, which is an e_mux
  assign p60_full_60 = ((read & !write) == 0)? full_59 :
    full_61;

  //control_reg_60, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_60 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_60 <= 0;
          else 
            full_60 <= p60_full_60;
    end


  //data_59, which is an e_mux
  assign p59_stage_59 = ((full_60 & ~clear_fifo) == 0)? data_in :
    stage_60;

  //data_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_59 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_59))
          if (sync_reset & full_59 & !((full_60 == 0) & read & write))
              stage_59 <= 0;
          else 
            stage_59 <= p59_stage_59;
    end


  //control_59, which is an e_mux
  assign p59_full_59 = ((read & !write) == 0)? full_58 :
    full_60;

  //control_reg_59, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_59 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_59 <= 0;
          else 
            full_59 <= p59_full_59;
    end


  //data_58, which is an e_mux
  assign p58_stage_58 = ((full_59 & ~clear_fifo) == 0)? data_in :
    stage_59;

  //data_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_58 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_58))
          if (sync_reset & full_58 & !((full_59 == 0) & read & write))
              stage_58 <= 0;
          else 
            stage_58 <= p58_stage_58;
    end


  //control_58, which is an e_mux
  assign p58_full_58 = ((read & !write) == 0)? full_57 :
    full_59;

  //control_reg_58, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_58 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_58 <= 0;
          else 
            full_58 <= p58_full_58;
    end


  //data_57, which is an e_mux
  assign p57_stage_57 = ((full_58 & ~clear_fifo) == 0)? data_in :
    stage_58;

  //data_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_57 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_57))
          if (sync_reset & full_57 & !((full_58 == 0) & read & write))
              stage_57 <= 0;
          else 
            stage_57 <= p57_stage_57;
    end


  //control_57, which is an e_mux
  assign p57_full_57 = ((read & !write) == 0)? full_56 :
    full_58;

  //control_reg_57, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_57 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_57 <= 0;
          else 
            full_57 <= p57_full_57;
    end


  //data_56, which is an e_mux
  assign p56_stage_56 = ((full_57 & ~clear_fifo) == 0)? data_in :
    stage_57;

  //data_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_56 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_56))
          if (sync_reset & full_56 & !((full_57 == 0) & read & write))
              stage_56 <= 0;
          else 
            stage_56 <= p56_stage_56;
    end


  //control_56, which is an e_mux
  assign p56_full_56 = ((read & !write) == 0)? full_55 :
    full_57;

  //control_reg_56, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_56 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_56 <= 0;
          else 
            full_56 <= p56_full_56;
    end


  //data_55, which is an e_mux
  assign p55_stage_55 = ((full_56 & ~clear_fifo) == 0)? data_in :
    stage_56;

  //data_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_55 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_55))
          if (sync_reset & full_55 & !((full_56 == 0) & read & write))
              stage_55 <= 0;
          else 
            stage_55 <= p55_stage_55;
    end


  //control_55, which is an e_mux
  assign p55_full_55 = ((read & !write) == 0)? full_54 :
    full_56;

  //control_reg_55, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_55 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_55 <= 0;
          else 
            full_55 <= p55_full_55;
    end


  //data_54, which is an e_mux
  assign p54_stage_54 = ((full_55 & ~clear_fifo) == 0)? data_in :
    stage_55;

  //data_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_54 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_54))
          if (sync_reset & full_54 & !((full_55 == 0) & read & write))
              stage_54 <= 0;
          else 
            stage_54 <= p54_stage_54;
    end


  //control_54, which is an e_mux
  assign p54_full_54 = ((read & !write) == 0)? full_53 :
    full_55;

  //control_reg_54, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_54 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_54 <= 0;
          else 
            full_54 <= p54_full_54;
    end


  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    stage_54;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    full_54;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_s1_arbitrator (
                                      // inputs:
                                       Medipix_sopc_burst_4_downstream_address_to_slave,
                                       Medipix_sopc_burst_4_downstream_arbitrationshare,
                                       Medipix_sopc_burst_4_downstream_burstcount,
                                       Medipix_sopc_burst_4_downstream_byteenable,
                                       Medipix_sopc_burst_4_downstream_latency_counter,
                                       Medipix_sopc_burst_4_downstream_nativeaddress,
                                       Medipix_sopc_burst_4_downstream_read,
                                       Medipix_sopc_burst_4_downstream_write,
                                       Medipix_sopc_burst_4_downstream_writedata,
                                       Medipix_sopc_burst_5_downstream_address_to_slave,
                                       Medipix_sopc_burst_5_downstream_arbitrationshare,
                                       Medipix_sopc_burst_5_downstream_burstcount,
                                       Medipix_sopc_burst_5_downstream_byteenable,
                                       Medipix_sopc_burst_5_downstream_latency_counter,
                                       Medipix_sopc_burst_5_downstream_nativeaddress,
                                       Medipix_sopc_burst_5_downstream_read,
                                       Medipix_sopc_burst_5_downstream_write,
                                       Medipix_sopc_burst_5_downstream_writedata,
                                       clk,
                                       clock_crossing_s1_endofpacket,
                                       clock_crossing_s1_readdata,
                                       clock_crossing_s1_readdatavalid,
                                       clock_crossing_s1_waitrequest,
                                       igor_mac_rx_master_address_to_slave,
                                       igor_mac_rx_master_byteenable,
                                       igor_mac_rx_master_write,
                                       igor_mac_rx_master_writedata,
                                       igor_mac_tx_master_address_to_slave,
                                       igor_mac_tx_master_latency_counter,
                                       igor_mac_tx_master_read,
                                       reset_n,

                                      // outputs:
                                       Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1,
                                       Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1,
                                       Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1,
                                       Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register,
                                       Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1,
                                       Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1,
                                       Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1,
                                       Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1,
                                       Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register,
                                       Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1,
                                       clock_crossing_s1_address,
                                       clock_crossing_s1_byteenable,
                                       clock_crossing_s1_endofpacket_from_sa,
                                       clock_crossing_s1_nativeaddress,
                                       clock_crossing_s1_read,
                                       clock_crossing_s1_readdata_from_sa,
                                       clock_crossing_s1_reset_n,
                                       clock_crossing_s1_waitrequest_from_sa,
                                       clock_crossing_s1_write,
                                       clock_crossing_s1_writedata,
                                       d1_clock_crossing_s1_end_xfer,
                                       igor_mac_rx_master_granted_clock_crossing_s1,
                                       igor_mac_rx_master_qualified_request_clock_crossing_s1,
                                       igor_mac_rx_master_requests_clock_crossing_s1,
                                       igor_mac_tx_master_granted_clock_crossing_s1,
                                       igor_mac_tx_master_qualified_request_clock_crossing_s1,
                                       igor_mac_tx_master_read_data_valid_clock_crossing_s1,
                                       igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register,
                                       igor_mac_tx_master_requests_clock_crossing_s1
                                    )
;

  output           Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1;
  output           Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1;
  output           Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1;
  output           Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register;
  output           Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1;
  output           Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1;
  output           Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1;
  output           Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1;
  output           Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register;
  output           Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1;
  output  [ 24: 0] clock_crossing_s1_address;
  output  [  3: 0] clock_crossing_s1_byteenable;
  output           clock_crossing_s1_endofpacket_from_sa;
  output  [ 24: 0] clock_crossing_s1_nativeaddress;
  output           clock_crossing_s1_read;
  output  [ 31: 0] clock_crossing_s1_readdata_from_sa;
  output           clock_crossing_s1_reset_n;
  output           clock_crossing_s1_waitrequest_from_sa;
  output           clock_crossing_s1_write;
  output  [ 31: 0] clock_crossing_s1_writedata;
  output           d1_clock_crossing_s1_end_xfer;
  output           igor_mac_rx_master_granted_clock_crossing_s1;
  output           igor_mac_rx_master_qualified_request_clock_crossing_s1;
  output           igor_mac_rx_master_requests_clock_crossing_s1;
  output           igor_mac_tx_master_granted_clock_crossing_s1;
  output           igor_mac_tx_master_qualified_request_clock_crossing_s1;
  output           igor_mac_tx_master_read_data_valid_clock_crossing_s1;
  output           igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register;
  output           igor_mac_tx_master_requests_clock_crossing_s1;
  input   [ 26: 0] Medipix_sopc_burst_4_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_4_downstream_arbitrationshare;
  input            Medipix_sopc_burst_4_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_4_downstream_byteenable;
  input            Medipix_sopc_burst_4_downstream_latency_counter;
  input   [ 26: 0] Medipix_sopc_burst_4_downstream_nativeaddress;
  input            Medipix_sopc_burst_4_downstream_read;
  input            Medipix_sopc_burst_4_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_4_downstream_writedata;
  input   [ 26: 0] Medipix_sopc_burst_5_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_5_downstream_arbitrationshare;
  input            Medipix_sopc_burst_5_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_5_downstream_byteenable;
  input            Medipix_sopc_burst_5_downstream_latency_counter;
  input   [ 26: 0] Medipix_sopc_burst_5_downstream_nativeaddress;
  input            Medipix_sopc_burst_5_downstream_read;
  input            Medipix_sopc_burst_5_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_5_downstream_writedata;
  input            clk;
  input            clock_crossing_s1_endofpacket;
  input   [ 31: 0] clock_crossing_s1_readdata;
  input            clock_crossing_s1_readdatavalid;
  input            clock_crossing_s1_waitrequest;
  input   [ 31: 0] igor_mac_rx_master_address_to_slave;
  input   [  3: 0] igor_mac_rx_master_byteenable;
  input            igor_mac_rx_master_write;
  input   [ 31: 0] igor_mac_rx_master_writedata;
  input   [ 31: 0] igor_mac_tx_master_address_to_slave;
  input            igor_mac_tx_master_latency_counter;
  input            igor_mac_tx_master_read;
  input            reset_n;

  wire             Medipix_sopc_burst_4_downstream_arbiterlock;
  wire             Medipix_sopc_burst_4_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_4_downstream_continuerequest;
  wire             Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_rdv_fifo_empty_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_rdv_fifo_output_from_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register;
  wire             Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_arbiterlock;
  wire             Medipix_sopc_burst_5_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_5_downstream_continuerequest;
  wire             Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_rdv_fifo_empty_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_rdv_fifo_output_from_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register;
  wire             Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1;
  wire    [ 24: 0] clock_crossing_s1_address;
  wire             clock_crossing_s1_allgrants;
  wire             clock_crossing_s1_allow_new_arb_cycle;
  wire             clock_crossing_s1_any_bursting_master_saved_grant;
  wire             clock_crossing_s1_any_continuerequest;
  reg     [  3: 0] clock_crossing_s1_arb_addend;
  wire             clock_crossing_s1_arb_counter_enable;
  reg     [  3: 0] clock_crossing_s1_arb_share_counter;
  wire    [  3: 0] clock_crossing_s1_arb_share_counter_next_value;
  wire    [  3: 0] clock_crossing_s1_arb_share_set_values;
  wire    [  3: 0] clock_crossing_s1_arb_winner;
  wire             clock_crossing_s1_arbitration_holdoff_internal;
  wire             clock_crossing_s1_beginbursttransfer_internal;
  wire             clock_crossing_s1_begins_xfer;
  wire    [  3: 0] clock_crossing_s1_byteenable;
  wire    [  7: 0] clock_crossing_s1_chosen_master_double_vector;
  wire    [  3: 0] clock_crossing_s1_chosen_master_rot_left;
  wire             clock_crossing_s1_end_xfer;
  wire             clock_crossing_s1_endofpacket_from_sa;
  wire             clock_crossing_s1_firsttransfer;
  wire    [  3: 0] clock_crossing_s1_grant_vector;
  wire             clock_crossing_s1_in_a_read_cycle;
  wire             clock_crossing_s1_in_a_write_cycle;
  wire    [  3: 0] clock_crossing_s1_master_qreq_vector;
  wire             clock_crossing_s1_move_on_to_next_transaction;
  wire    [ 24: 0] clock_crossing_s1_nativeaddress;
  wire             clock_crossing_s1_non_bursting_master_requests;
  wire             clock_crossing_s1_read;
  wire    [ 31: 0] clock_crossing_s1_readdata_from_sa;
  wire             clock_crossing_s1_readdatavalid_from_sa;
  reg              clock_crossing_s1_reg_firsttransfer;
  wire             clock_crossing_s1_reset_n;
  reg     [  3: 0] clock_crossing_s1_saved_chosen_master_vector;
  reg              clock_crossing_s1_slavearbiterlockenable;
  wire             clock_crossing_s1_slavearbiterlockenable2;
  wire             clock_crossing_s1_unreg_firsttransfer;
  wire             clock_crossing_s1_waitrequest_from_sa;
  wire             clock_crossing_s1_waits_for_read;
  wire             clock_crossing_s1_waits_for_write;
  wire             clock_crossing_s1_write;
  wire    [ 31: 0] clock_crossing_s1_writedata;
  reg              d1_clock_crossing_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_clock_crossing_s1;
  wire             igor_mac_rx_master_arbiterlock;
  wire             igor_mac_rx_master_arbiterlock2;
  wire             igor_mac_rx_master_continuerequest;
  wire             igor_mac_rx_master_granted_clock_crossing_s1;
  wire             igor_mac_rx_master_qualified_request_clock_crossing_s1;
  wire             igor_mac_rx_master_requests_clock_crossing_s1;
  wire             igor_mac_rx_master_saved_grant_clock_crossing_s1;
  wire             igor_mac_tx_master_arbiterlock;
  wire             igor_mac_tx_master_arbiterlock2;
  wire             igor_mac_tx_master_continuerequest;
  wire             igor_mac_tx_master_granted_clock_crossing_s1;
  wire             igor_mac_tx_master_qualified_request_clock_crossing_s1;
  wire             igor_mac_tx_master_rdv_fifo_empty_clock_crossing_s1;
  wire             igor_mac_tx_master_rdv_fifo_output_from_clock_crossing_s1;
  wire             igor_mac_tx_master_read_data_valid_clock_crossing_s1;
  wire             igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register;
  wire             igor_mac_tx_master_requests_clock_crossing_s1;
  wire             igor_mac_tx_master_saved_grant_clock_crossing_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1;
  reg              last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1;
  reg              last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1;
  reg              last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1;
  wire    [ 26: 0] shifted_address_to_clock_crossing_s1_from_Medipix_sopc_burst_4_downstream;
  wire    [ 26: 0] shifted_address_to_clock_crossing_s1_from_Medipix_sopc_burst_5_downstream;
  wire    [ 31: 0] shifted_address_to_clock_crossing_s1_from_igor_mac_rx_master;
  wire    [ 31: 0] shifted_address_to_clock_crossing_s1_from_igor_mac_tx_master;
  wire             wait_for_clock_crossing_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~clock_crossing_s1_end_xfer;
    end


  assign clock_crossing_s1_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1 | Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1 | igor_mac_rx_master_qualified_request_clock_crossing_s1 | igor_mac_tx_master_qualified_request_clock_crossing_s1));
  //assign clock_crossing_s1_readdata_from_sa = clock_crossing_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_s1_readdata_from_sa = clock_crossing_s1_readdata;

  assign Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1 = (1) & (Medipix_sopc_burst_4_downstream_read | Medipix_sopc_burst_4_downstream_write);
  //assign clock_crossing_s1_waitrequest_from_sa = clock_crossing_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_s1_waitrequest_from_sa = clock_crossing_s1_waitrequest;

  //assign clock_crossing_s1_readdatavalid_from_sa = clock_crossing_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_s1_readdatavalid_from_sa = clock_crossing_s1_readdatavalid;

  //clock_crossing_s1_arb_share_counter set values, which is an e_mux
  assign clock_crossing_s1_arb_share_set_values = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_arbitrationshare :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_arbitrationshare :
    (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_arbitrationshare :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_arbitrationshare :
    (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_arbitrationshare :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_arbitrationshare :
    (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_arbitrationshare :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_arbitrationshare :
    1;

  //clock_crossing_s1_non_bursting_master_requests mux, which is an e_mux
  assign clock_crossing_s1_non_bursting_master_requests = 0 |
    igor_mac_rx_master_requests_clock_crossing_s1 |
    igor_mac_tx_master_requests_clock_crossing_s1 |
    igor_mac_rx_master_requests_clock_crossing_s1 |
    igor_mac_tx_master_requests_clock_crossing_s1 |
    igor_mac_rx_master_requests_clock_crossing_s1 |
    igor_mac_tx_master_requests_clock_crossing_s1 |
    igor_mac_rx_master_requests_clock_crossing_s1 |
    igor_mac_tx_master_requests_clock_crossing_s1;

  //clock_crossing_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign clock_crossing_s1_any_bursting_master_saved_grant = Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 |
    Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1;

  //clock_crossing_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign clock_crossing_s1_arb_share_counter_next_value = clock_crossing_s1_firsttransfer ? (clock_crossing_s1_arb_share_set_values - 1) : |clock_crossing_s1_arb_share_counter ? (clock_crossing_s1_arb_share_counter - 1) : 0;

  //clock_crossing_s1_allgrants all slave grants, which is an e_mux
  assign clock_crossing_s1_allgrants = (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector) |
    (|clock_crossing_s1_grant_vector);

  //clock_crossing_s1_end_xfer assignment, which is an e_assign
  assign clock_crossing_s1_end_xfer = ~(clock_crossing_s1_waits_for_read | clock_crossing_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_clock_crossing_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_clock_crossing_s1 = clock_crossing_s1_end_xfer & (~clock_crossing_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //clock_crossing_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign clock_crossing_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_clock_crossing_s1 & clock_crossing_s1_allgrants) | (end_xfer_arb_share_counter_term_clock_crossing_s1 & ~clock_crossing_s1_non_bursting_master_requests);

  //clock_crossing_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_s1_arb_share_counter <= 0;
      else if (clock_crossing_s1_arb_counter_enable)
          clock_crossing_s1_arb_share_counter <= clock_crossing_s1_arb_share_counter_next_value;
    end


  //clock_crossing_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_s1_slavearbiterlockenable <= 0;
      else if ((|clock_crossing_s1_master_qreq_vector & end_xfer_arb_share_counter_term_clock_crossing_s1) | (end_xfer_arb_share_counter_term_clock_crossing_s1 & ~clock_crossing_s1_non_bursting_master_requests))
          clock_crossing_s1_slavearbiterlockenable <= |clock_crossing_s1_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_4/downstream clock_crossing/s1 arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_arbiterlock = clock_crossing_s1_slavearbiterlockenable & Medipix_sopc_burst_4_downstream_continuerequest;

  //clock_crossing_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign clock_crossing_s1_slavearbiterlockenable2 = |clock_crossing_s1_arb_share_counter_next_value;

  //Medipix_sopc_burst_4/downstream clock_crossing/s1 arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_arbiterlock2 = clock_crossing_s1_slavearbiterlockenable2 & Medipix_sopc_burst_4_downstream_continuerequest;

  //Medipix_sopc_burst_5/downstream clock_crossing/s1 arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_arbiterlock = clock_crossing_s1_slavearbiterlockenable & Medipix_sopc_burst_5_downstream_continuerequest;

  //Medipix_sopc_burst_5/downstream clock_crossing/s1 arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_arbiterlock2 = clock_crossing_s1_slavearbiterlockenable2 & Medipix_sopc_burst_5_downstream_continuerequest;

  //Medipix_sopc_burst_5/downstream granted clock_crossing/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1 <= 0;
      else 
        last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1 <= Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1 ? 1 : (clock_crossing_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1;
    end


  //Medipix_sopc_burst_5_downstream_continuerequest continued request, which is an e_mux
  assign Medipix_sopc_burst_5_downstream_continuerequest = (last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1 & 1) |
    (last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1 & 1) |
    (last_cycle_Medipix_sopc_burst_5_downstream_granted_slave_clock_crossing_s1 & 1);

  //clock_crossing_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign clock_crossing_s1_any_continuerequest = Medipix_sopc_burst_5_downstream_continuerequest |
    igor_mac_rx_master_continuerequest |
    igor_mac_tx_master_continuerequest |
    Medipix_sopc_burst_4_downstream_continuerequest |
    igor_mac_rx_master_continuerequest |
    igor_mac_tx_master_continuerequest |
    Medipix_sopc_burst_4_downstream_continuerequest |
    Medipix_sopc_burst_5_downstream_continuerequest |
    igor_mac_tx_master_continuerequest |
    Medipix_sopc_burst_4_downstream_continuerequest |
    Medipix_sopc_burst_5_downstream_continuerequest |
    igor_mac_rx_master_continuerequest;

  //igor_mac/rx_master clock_crossing/s1 arbiterlock, which is an e_assign
  assign igor_mac_rx_master_arbiterlock = clock_crossing_s1_slavearbiterlockenable & igor_mac_rx_master_continuerequest;

  //igor_mac/rx_master clock_crossing/s1 arbiterlock2, which is an e_assign
  assign igor_mac_rx_master_arbiterlock2 = clock_crossing_s1_slavearbiterlockenable2 & igor_mac_rx_master_continuerequest;

  //igor_mac/rx_master granted clock_crossing/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1 <= 0;
      else 
        last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1 <= igor_mac_rx_master_saved_grant_clock_crossing_s1 ? 1 : (clock_crossing_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1;
    end


  //igor_mac_rx_master_continuerequest continued request, which is an e_mux
  assign igor_mac_rx_master_continuerequest = (last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1 & igor_mac_rx_master_requests_clock_crossing_s1) |
    (last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1 & igor_mac_rx_master_requests_clock_crossing_s1) |
    (last_cycle_igor_mac_rx_master_granted_slave_clock_crossing_s1 & igor_mac_rx_master_requests_clock_crossing_s1);

  //igor_mac/tx_master clock_crossing/s1 arbiterlock, which is an e_assign
  assign igor_mac_tx_master_arbiterlock = clock_crossing_s1_slavearbiterlockenable & igor_mac_tx_master_continuerequest;

  //igor_mac/tx_master clock_crossing/s1 arbiterlock2, which is an e_assign
  assign igor_mac_tx_master_arbiterlock2 = clock_crossing_s1_slavearbiterlockenable2 & igor_mac_tx_master_continuerequest;

  //igor_mac/tx_master granted clock_crossing/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1 <= 0;
      else 
        last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1 <= igor_mac_tx_master_saved_grant_clock_crossing_s1 ? 1 : (clock_crossing_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1;
    end


  //igor_mac_tx_master_continuerequest continued request, which is an e_mux
  assign igor_mac_tx_master_continuerequest = (last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1 & igor_mac_tx_master_requests_clock_crossing_s1) |
    (last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1 & igor_mac_tx_master_requests_clock_crossing_s1) |
    (last_cycle_igor_mac_tx_master_granted_slave_clock_crossing_s1 & igor_mac_tx_master_requests_clock_crossing_s1);

  assign Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1 = Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1 & ~((Medipix_sopc_burst_4_downstream_read & ((Medipix_sopc_burst_4_downstream_latency_counter != 0) | (1 < Medipix_sopc_burst_4_downstream_latency_counter))) | Medipix_sopc_burst_5_downstream_arbiterlock | igor_mac_rx_master_arbiterlock | igor_mac_tx_master_arbiterlock);
  //unique name for clock_crossing_s1_move_on_to_next_transaction, which is an e_assign
  assign clock_crossing_s1_move_on_to_next_transaction = clock_crossing_s1_readdatavalid_from_sa;

  //rdv_fifo_for_Medipix_sopc_burst_4_downstream_to_clock_crossing_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_Medipix_sopc_burst_4_downstream_to_clock_crossing_s1_module rdv_fifo_for_Medipix_sopc_burst_4_downstream_to_clock_crossing_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1),
      .data_out             (Medipix_sopc_burst_4_downstream_rdv_fifo_output_from_clock_crossing_s1),
      .empty                (),
      .fifo_contains_ones_n (Medipix_sopc_burst_4_downstream_rdv_fifo_empty_clock_crossing_s1),
      .full                 (),
      .read                 (clock_crossing_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_s1_waits_for_read)
    );

  assign Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register = ~Medipix_sopc_burst_4_downstream_rdv_fifo_empty_clock_crossing_s1;
  //local readdatavalid Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1, which is an e_mux
  assign Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1 = (clock_crossing_s1_readdatavalid_from_sa & Medipix_sopc_burst_4_downstream_rdv_fifo_output_from_clock_crossing_s1) & ~ Medipix_sopc_burst_4_downstream_rdv_fifo_empty_clock_crossing_s1;

  //clock_crossing_s1_writedata mux, which is an e_mux
  assign clock_crossing_s1_writedata = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_writedata :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_writedata :
    igor_mac_rx_master_writedata;

  //assign clock_crossing_s1_endofpacket_from_sa = clock_crossing_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_s1_endofpacket_from_sa = clock_crossing_s1_endofpacket;

  assign Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1 = (1) & (Medipix_sopc_burst_5_downstream_read | Medipix_sopc_burst_5_downstream_write);
  //Medipix_sopc_burst_4/downstream granted clock_crossing/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1 <= 0;
      else 
        last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1 <= Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 ? 1 : (clock_crossing_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1;
    end


  //Medipix_sopc_burst_4_downstream_continuerequest continued request, which is an e_mux
  assign Medipix_sopc_burst_4_downstream_continuerequest = (last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1 & 1) |
    (last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1 & 1) |
    (last_cycle_Medipix_sopc_burst_4_downstream_granted_slave_clock_crossing_s1 & 1);

  assign Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1 = Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1 & ~((Medipix_sopc_burst_5_downstream_read & ((Medipix_sopc_burst_5_downstream_latency_counter != 0) | (1 < Medipix_sopc_burst_5_downstream_latency_counter))) | Medipix_sopc_burst_4_downstream_arbiterlock | igor_mac_rx_master_arbiterlock | igor_mac_tx_master_arbiterlock);
  //rdv_fifo_for_Medipix_sopc_burst_5_downstream_to_clock_crossing_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_Medipix_sopc_burst_5_downstream_to_clock_crossing_s1_module rdv_fifo_for_Medipix_sopc_burst_5_downstream_to_clock_crossing_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1),
      .data_out             (Medipix_sopc_burst_5_downstream_rdv_fifo_output_from_clock_crossing_s1),
      .empty                (),
      .fifo_contains_ones_n (Medipix_sopc_burst_5_downstream_rdv_fifo_empty_clock_crossing_s1),
      .full                 (),
      .read                 (clock_crossing_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_s1_waits_for_read)
    );

  assign Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register = ~Medipix_sopc_burst_5_downstream_rdv_fifo_empty_clock_crossing_s1;
  //local readdatavalid Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1, which is an e_mux
  assign Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1 = (clock_crossing_s1_readdatavalid_from_sa & Medipix_sopc_burst_5_downstream_rdv_fifo_output_from_clock_crossing_s1) & ~ Medipix_sopc_burst_5_downstream_rdv_fifo_empty_clock_crossing_s1;

  assign igor_mac_rx_master_requests_clock_crossing_s1 = (({igor_mac_rx_master_address_to_slave[31 : 27] , 27'b0} == 32'h0) & (igor_mac_rx_master_write)) & igor_mac_rx_master_write;
  assign igor_mac_rx_master_qualified_request_clock_crossing_s1 = igor_mac_rx_master_requests_clock_crossing_s1 & ~(Medipix_sopc_burst_4_downstream_arbiterlock | Medipix_sopc_burst_5_downstream_arbiterlock | igor_mac_tx_master_arbiterlock);
  assign igor_mac_tx_master_requests_clock_crossing_s1 = (({igor_mac_tx_master_address_to_slave[31 : 27] , 27'b0} == 32'h0) & (igor_mac_tx_master_read)) & igor_mac_tx_master_read;
  assign igor_mac_tx_master_qualified_request_clock_crossing_s1 = igor_mac_tx_master_requests_clock_crossing_s1 & ~((igor_mac_tx_master_read & ((igor_mac_tx_master_latency_counter != 0) | (1 < igor_mac_tx_master_latency_counter))) | Medipix_sopc_burst_4_downstream_arbiterlock | Medipix_sopc_burst_5_downstream_arbiterlock | igor_mac_rx_master_arbiterlock);
  //rdv_fifo_for_igor_mac_tx_master_to_clock_crossing_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_igor_mac_tx_master_to_clock_crossing_s1_module rdv_fifo_for_igor_mac_tx_master_to_clock_crossing_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (igor_mac_tx_master_granted_clock_crossing_s1),
      .data_out             (igor_mac_tx_master_rdv_fifo_output_from_clock_crossing_s1),
      .empty                (),
      .fifo_contains_ones_n (igor_mac_tx_master_rdv_fifo_empty_clock_crossing_s1),
      .full                 (),
      .read                 (clock_crossing_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_s1_waits_for_read)
    );

  assign igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register = ~igor_mac_tx_master_rdv_fifo_empty_clock_crossing_s1;
  //local readdatavalid igor_mac_tx_master_read_data_valid_clock_crossing_s1, which is an e_mux
  assign igor_mac_tx_master_read_data_valid_clock_crossing_s1 = (clock_crossing_s1_readdatavalid_from_sa & igor_mac_tx_master_rdv_fifo_output_from_clock_crossing_s1) & ~ igor_mac_tx_master_rdv_fifo_empty_clock_crossing_s1;

  //allow new arb cycle for clock_crossing/s1, which is an e_assign
  assign clock_crossing_s1_allow_new_arb_cycle = ~Medipix_sopc_burst_4_downstream_arbiterlock & ~Medipix_sopc_burst_5_downstream_arbiterlock & ~igor_mac_rx_master_arbiterlock & ~igor_mac_tx_master_arbiterlock;

  //igor_mac/tx_master assignment into master qualified-requests vector for clock_crossing/s1, which is an e_assign
  assign clock_crossing_s1_master_qreq_vector[0] = igor_mac_tx_master_qualified_request_clock_crossing_s1;

  //igor_mac/tx_master grant clock_crossing/s1, which is an e_assign
  assign igor_mac_tx_master_granted_clock_crossing_s1 = clock_crossing_s1_grant_vector[0];

  //igor_mac/tx_master saved-grant clock_crossing/s1, which is an e_assign
  assign igor_mac_tx_master_saved_grant_clock_crossing_s1 = clock_crossing_s1_arb_winner[0] && igor_mac_tx_master_requests_clock_crossing_s1;

  //igor_mac/rx_master assignment into master qualified-requests vector for clock_crossing/s1, which is an e_assign
  assign clock_crossing_s1_master_qreq_vector[1] = igor_mac_rx_master_qualified_request_clock_crossing_s1;

  //igor_mac/rx_master grant clock_crossing/s1, which is an e_assign
  assign igor_mac_rx_master_granted_clock_crossing_s1 = clock_crossing_s1_grant_vector[1];

  //igor_mac/rx_master saved-grant clock_crossing/s1, which is an e_assign
  assign igor_mac_rx_master_saved_grant_clock_crossing_s1 = clock_crossing_s1_arb_winner[1] && igor_mac_rx_master_requests_clock_crossing_s1;

  //Medipix_sopc_burst_5/downstream assignment into master qualified-requests vector for clock_crossing/s1, which is an e_assign
  assign clock_crossing_s1_master_qreq_vector[2] = Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1;

  //Medipix_sopc_burst_5/downstream grant clock_crossing/s1, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 = clock_crossing_s1_grant_vector[2];

  //Medipix_sopc_burst_5/downstream saved-grant clock_crossing/s1, which is an e_assign
  assign Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1 = clock_crossing_s1_arb_winner[2];

  //Medipix_sopc_burst_4/downstream assignment into master qualified-requests vector for clock_crossing/s1, which is an e_assign
  assign clock_crossing_s1_master_qreq_vector[3] = Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1;

  //Medipix_sopc_burst_4/downstream grant clock_crossing/s1, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 = clock_crossing_s1_grant_vector[3];

  //Medipix_sopc_burst_4/downstream saved-grant clock_crossing/s1, which is an e_assign
  assign Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 = clock_crossing_s1_arb_winner[3];

  //clock_crossing/s1 chosen-master double-vector, which is an e_assign
  assign clock_crossing_s1_chosen_master_double_vector = {clock_crossing_s1_master_qreq_vector, clock_crossing_s1_master_qreq_vector} & ({~clock_crossing_s1_master_qreq_vector, ~clock_crossing_s1_master_qreq_vector} + clock_crossing_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign clock_crossing_s1_arb_winner = (clock_crossing_s1_allow_new_arb_cycle & | clock_crossing_s1_grant_vector) ? clock_crossing_s1_grant_vector : clock_crossing_s1_saved_chosen_master_vector;

  //saved clock_crossing_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_s1_saved_chosen_master_vector <= 0;
      else if (clock_crossing_s1_allow_new_arb_cycle)
          clock_crossing_s1_saved_chosen_master_vector <= |clock_crossing_s1_grant_vector ? clock_crossing_s1_grant_vector : clock_crossing_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign clock_crossing_s1_grant_vector = {(clock_crossing_s1_chosen_master_double_vector[3] | clock_crossing_s1_chosen_master_double_vector[7]),
    (clock_crossing_s1_chosen_master_double_vector[2] | clock_crossing_s1_chosen_master_double_vector[6]),
    (clock_crossing_s1_chosen_master_double_vector[1] | clock_crossing_s1_chosen_master_double_vector[5]),
    (clock_crossing_s1_chosen_master_double_vector[0] | clock_crossing_s1_chosen_master_double_vector[4])};

  //clock_crossing/s1 chosen master rotated left, which is an e_assign
  assign clock_crossing_s1_chosen_master_rot_left = (clock_crossing_s1_arb_winner << 1) ? (clock_crossing_s1_arb_winner << 1) : 1;

  //clock_crossing/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_s1_arb_addend <= 1;
      else if (|clock_crossing_s1_grant_vector)
          clock_crossing_s1_arb_addend <= clock_crossing_s1_end_xfer? clock_crossing_s1_chosen_master_rot_left : clock_crossing_s1_grant_vector;
    end


  //clock_crossing_s1_reset_n assignment, which is an e_assign
  assign clock_crossing_s1_reset_n = reset_n;

  //clock_crossing_s1_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_s1_firsttransfer = clock_crossing_s1_begins_xfer ? clock_crossing_s1_unreg_firsttransfer : clock_crossing_s1_reg_firsttransfer;

  //clock_crossing_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_s1_unreg_firsttransfer = ~(clock_crossing_s1_slavearbiterlockenable & clock_crossing_s1_any_continuerequest);

  //clock_crossing_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_s1_reg_firsttransfer <= 1'b1;
      else if (clock_crossing_s1_begins_xfer)
          clock_crossing_s1_reg_firsttransfer <= clock_crossing_s1_unreg_firsttransfer;
    end


  //clock_crossing_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign clock_crossing_s1_beginbursttransfer_internal = clock_crossing_s1_begins_xfer;

  //clock_crossing_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign clock_crossing_s1_arbitration_holdoff_internal = clock_crossing_s1_begins_xfer & clock_crossing_s1_firsttransfer;

  //clock_crossing_s1_read assignment, which is an e_mux
  assign clock_crossing_s1_read = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_4_downstream_read) | (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_5_downstream_read) | (igor_mac_tx_master_granted_clock_crossing_s1 & igor_mac_tx_master_read);

  //clock_crossing_s1_write assignment, which is an e_mux
  assign clock_crossing_s1_write = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_4_downstream_write) | (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_5_downstream_write) | (igor_mac_rx_master_granted_clock_crossing_s1 & igor_mac_rx_master_write);

  assign shifted_address_to_clock_crossing_s1_from_Medipix_sopc_burst_4_downstream = Medipix_sopc_burst_4_downstream_address_to_slave;
  //clock_crossing_s1_address mux, which is an e_mux
  assign clock_crossing_s1_address = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? (shifted_address_to_clock_crossing_s1_from_Medipix_sopc_burst_4_downstream >> 2) :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? (shifted_address_to_clock_crossing_s1_from_Medipix_sopc_burst_5_downstream >> 2) :
    (igor_mac_rx_master_granted_clock_crossing_s1)? (shifted_address_to_clock_crossing_s1_from_igor_mac_rx_master >> 2) :
    (shifted_address_to_clock_crossing_s1_from_igor_mac_tx_master >> 2);

  assign shifted_address_to_clock_crossing_s1_from_Medipix_sopc_burst_5_downstream = Medipix_sopc_burst_5_downstream_address_to_slave;
  assign shifted_address_to_clock_crossing_s1_from_igor_mac_rx_master = igor_mac_rx_master_address_to_slave;
  assign shifted_address_to_clock_crossing_s1_from_igor_mac_tx_master = igor_mac_tx_master_address_to_slave;
  //slaveid clock_crossing_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign clock_crossing_s1_nativeaddress = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_nativeaddress :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_nativeaddress :
    (igor_mac_rx_master_granted_clock_crossing_s1)? (igor_mac_rx_master_address_to_slave >> 2) :
    (igor_mac_tx_master_address_to_slave >> 2);

  //d1_clock_crossing_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_clock_crossing_s1_end_xfer <= 1;
      else 
        d1_clock_crossing_s1_end_xfer <= clock_crossing_s1_end_xfer;
    end


  //clock_crossing_s1_waits_for_read in a cycle, which is an e_mux
  assign clock_crossing_s1_waits_for_read = clock_crossing_s1_in_a_read_cycle & clock_crossing_s1_waitrequest_from_sa;

  //clock_crossing_s1_in_a_read_cycle assignment, which is an e_assign
  assign clock_crossing_s1_in_a_read_cycle = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_4_downstream_read) | (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_5_downstream_read) | (igor_mac_tx_master_granted_clock_crossing_s1 & igor_mac_tx_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = clock_crossing_s1_in_a_read_cycle;

  //clock_crossing_s1_waits_for_write in a cycle, which is an e_mux
  assign clock_crossing_s1_waits_for_write = clock_crossing_s1_in_a_write_cycle & clock_crossing_s1_waitrequest_from_sa;

  //clock_crossing_s1_in_a_write_cycle assignment, which is an e_assign
  assign clock_crossing_s1_in_a_write_cycle = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_4_downstream_write) | (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 & Medipix_sopc_burst_5_downstream_write) | (igor_mac_rx_master_granted_clock_crossing_s1 & igor_mac_rx_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = clock_crossing_s1_in_a_write_cycle;

  assign wait_for_clock_crossing_s1_counter = 0;
  //clock_crossing_s1_byteenable byte enable port mux, which is an e_mux
  assign clock_crossing_s1_byteenable = (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_4_downstream_byteenable :
    (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1)? Medipix_sopc_burst_5_downstream_byteenable :
    (igor_mac_rx_master_granted_clock_crossing_s1)? igor_mac_rx_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_4/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1 && (Medipix_sopc_burst_4_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_4/downstream drove 0 on its 'arbitrationshare' port while accessing slave clock_crossing/s1", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_4/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1 && (Medipix_sopc_burst_4_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_4/downstream drove 0 on its 'burstcount' port while accessing slave clock_crossing/s1", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1 && (Medipix_sopc_burst_5_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_5/downstream drove 0 on its 'arbitrationshare' port while accessing slave clock_crossing/s1", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_5/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1 && (Medipix_sopc_burst_5_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_5/downstream drove 0 on its 'burstcount' port while accessing slave clock_crossing/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1 + Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1 + igor_mac_rx_master_granted_clock_crossing_s1 + igor_mac_tx_master_granted_clock_crossing_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_4_downstream_saved_grant_clock_crossing_s1 + Medipix_sopc_burst_5_downstream_saved_grant_clock_crossing_s1 + igor_mac_rx_master_saved_grant_clock_crossing_s1 + igor_mac_tx_master_saved_grant_clock_crossing_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_m1_arbitrator (
                                      // inputs:
                                       clk,
                                       clock_crossing_m1_address,
                                       clock_crossing_m1_byteenable,
                                       clock_crossing_m1_granted_ram_s1,
                                       clock_crossing_m1_qualified_request_ram_s1,
                                       clock_crossing_m1_read,
                                       clock_crossing_m1_read_data_valid_ram_s1,
                                       clock_crossing_m1_read_data_valid_ram_s1_shift_register,
                                       clock_crossing_m1_requests_ram_s1,
                                       clock_crossing_m1_write,
                                       clock_crossing_m1_writedata,
                                       d1_ram_s1_end_xfer,
                                       ram_s1_readdata_from_sa,
                                       ram_s1_waitrequest_n_from_sa,
                                       reset_n,

                                      // outputs:
                                       clock_crossing_m1_address_to_slave,
                                       clock_crossing_m1_latency_counter,
                                       clock_crossing_m1_readdata,
                                       clock_crossing_m1_readdatavalid,
                                       clock_crossing_m1_reset_n,
                                       clock_crossing_m1_waitrequest
                                    )
;

  output  [ 26: 0] clock_crossing_m1_address_to_slave;
  output           clock_crossing_m1_latency_counter;
  output  [ 31: 0] clock_crossing_m1_readdata;
  output           clock_crossing_m1_readdatavalid;
  output           clock_crossing_m1_reset_n;
  output           clock_crossing_m1_waitrequest;
  input            clk;
  input   [ 26: 0] clock_crossing_m1_address;
  input   [  3: 0] clock_crossing_m1_byteenable;
  input            clock_crossing_m1_granted_ram_s1;
  input            clock_crossing_m1_qualified_request_ram_s1;
  input            clock_crossing_m1_read;
  input            clock_crossing_m1_read_data_valid_ram_s1;
  input            clock_crossing_m1_read_data_valid_ram_s1_shift_register;
  input            clock_crossing_m1_requests_ram_s1;
  input            clock_crossing_m1_write;
  input   [ 31: 0] clock_crossing_m1_writedata;
  input            d1_ram_s1_end_xfer;
  input   [ 31: 0] ram_s1_readdata_from_sa;
  input            ram_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] clock_crossing_m1_address_last_time;
  wire    [ 26: 0] clock_crossing_m1_address_to_slave;
  reg     [  3: 0] clock_crossing_m1_byteenable_last_time;
  wire             clock_crossing_m1_latency_counter;
  reg              clock_crossing_m1_read_last_time;
  wire    [ 31: 0] clock_crossing_m1_readdata;
  wire             clock_crossing_m1_readdatavalid;
  wire             clock_crossing_m1_reset_n;
  wire             clock_crossing_m1_run;
  wire             clock_crossing_m1_waitrequest;
  reg              clock_crossing_m1_write_last_time;
  reg     [ 31: 0] clock_crossing_m1_writedata_last_time;
  wire             pre_flush_clock_crossing_m1_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (clock_crossing_m1_qualified_request_ram_s1 | ~clock_crossing_m1_requests_ram_s1) & ((~clock_crossing_m1_qualified_request_ram_s1 | ~(clock_crossing_m1_read | clock_crossing_m1_write) | (1 & ram_s1_waitrequest_n_from_sa & (clock_crossing_m1_read | clock_crossing_m1_write)))) & ((~clock_crossing_m1_qualified_request_ram_s1 | ~(clock_crossing_m1_read | clock_crossing_m1_write) | (1 & ram_s1_waitrequest_n_from_sa & (clock_crossing_m1_read | clock_crossing_m1_write))));

  //cascaded wait assignment, which is an e_assign
  assign clock_crossing_m1_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign clock_crossing_m1_address_to_slave = clock_crossing_m1_address[26 : 0];

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_clock_crossing_m1_readdatavalid = clock_crossing_m1_read_data_valid_ram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign clock_crossing_m1_readdatavalid = 0 |
    pre_flush_clock_crossing_m1_readdatavalid;

  //clock_crossing/m1 readdata mux, which is an e_mux
  assign clock_crossing_m1_readdata = ram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign clock_crossing_m1_waitrequest = ~clock_crossing_m1_run;

  //latent max counter, which is an e_assign
  assign clock_crossing_m1_latency_counter = 0;

  //clock_crossing_m1_reset_n assignment, which is an e_assign
  assign clock_crossing_m1_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_m1_address_last_time <= 0;
      else 
        clock_crossing_m1_address_last_time <= clock_crossing_m1_address;
    end


  //clock_crossing/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= clock_crossing_m1_waitrequest & (clock_crossing_m1_read | clock_crossing_m1_write);
    end


  //clock_crossing_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_m1_address != clock_crossing_m1_address_last_time))
        begin
          $write("%0d ns: clock_crossing_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_m1_byteenable_last_time <= 0;
      else 
        clock_crossing_m1_byteenable_last_time <= clock_crossing_m1_byteenable;
    end


  //clock_crossing_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_m1_byteenable != clock_crossing_m1_byteenable_last_time))
        begin
          $write("%0d ns: clock_crossing_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_m1_read_last_time <= 0;
      else 
        clock_crossing_m1_read_last_time <= clock_crossing_m1_read;
    end


  //clock_crossing_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_m1_read != clock_crossing_m1_read_last_time))
        begin
          $write("%0d ns: clock_crossing_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_m1_write_last_time <= 0;
      else 
        clock_crossing_m1_write_last_time <= clock_crossing_m1_write;
    end


  //clock_crossing_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_m1_write != clock_crossing_m1_write_last_time))
        begin
          $write("%0d ns: clock_crossing_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_m1_writedata_last_time <= 0;
      else 
        clock_crossing_m1_writedata_last_time <= clock_crossing_m1_writedata;
    end


  //clock_crossing_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_m1_writedata != clock_crossing_m1_writedata_last_time) & clock_crossing_m1_write)
        begin
          $write("%0d ns: clock_crossing_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_linux_jtag_debug_module_arbitrator (
                                                // inputs:
                                                 Medipix_sopc_burst_0_downstream_address_to_slave,
                                                 Medipix_sopc_burst_0_downstream_arbitrationshare,
                                                 Medipix_sopc_burst_0_downstream_burstcount,
                                                 Medipix_sopc_burst_0_downstream_byteenable,
                                                 Medipix_sopc_burst_0_downstream_debugaccess,
                                                 Medipix_sopc_burst_0_downstream_latency_counter,
                                                 Medipix_sopc_burst_0_downstream_read,
                                                 Medipix_sopc_burst_0_downstream_write,
                                                 Medipix_sopc_burst_0_downstream_writedata,
                                                 Medipix_sopc_burst_1_downstream_address_to_slave,
                                                 Medipix_sopc_burst_1_downstream_arbitrationshare,
                                                 Medipix_sopc_burst_1_downstream_burstcount,
                                                 Medipix_sopc_burst_1_downstream_byteenable,
                                                 Medipix_sopc_burst_1_downstream_debugaccess,
                                                 Medipix_sopc_burst_1_downstream_latency_counter,
                                                 Medipix_sopc_burst_1_downstream_read,
                                                 Medipix_sopc_burst_1_downstream_write,
                                                 Medipix_sopc_burst_1_downstream_writedata,
                                                 clk,
                                                 cpu_linux_jtag_debug_module_readdata,
                                                 cpu_linux_jtag_debug_module_resetrequest,
                                                 reset_n,

                                                // outputs:
                                                 Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module,
                                                 Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module,
                                                 cpu_linux_jtag_debug_module_address,
                                                 cpu_linux_jtag_debug_module_begintransfer,
                                                 cpu_linux_jtag_debug_module_byteenable,
                                                 cpu_linux_jtag_debug_module_chipselect,
                                                 cpu_linux_jtag_debug_module_debugaccess,
                                                 cpu_linux_jtag_debug_module_readdata_from_sa,
                                                 cpu_linux_jtag_debug_module_reset_n,
                                                 cpu_linux_jtag_debug_module_resetrequest_from_sa,
                                                 cpu_linux_jtag_debug_module_write,
                                                 cpu_linux_jtag_debug_module_writedata,
                                                 d1_cpu_linux_jtag_debug_module_end_xfer
                                              )
;

  output           Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  output           Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module;
  output  [  8: 0] cpu_linux_jtag_debug_module_address;
  output           cpu_linux_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_linux_jtag_debug_module_byteenable;
  output           cpu_linux_jtag_debug_module_chipselect;
  output           cpu_linux_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_linux_jtag_debug_module_readdata_from_sa;
  output           cpu_linux_jtag_debug_module_reset_n;
  output           cpu_linux_jtag_debug_module_resetrequest_from_sa;
  output           cpu_linux_jtag_debug_module_write;
  output  [ 31: 0] cpu_linux_jtag_debug_module_writedata;
  output           d1_cpu_linux_jtag_debug_module_end_xfer;
  input   [ 10: 0] Medipix_sopc_burst_0_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_0_downstream_arbitrationshare;
  input            Medipix_sopc_burst_0_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_0_downstream_byteenable;
  input            Medipix_sopc_burst_0_downstream_debugaccess;
  input            Medipix_sopc_burst_0_downstream_latency_counter;
  input            Medipix_sopc_burst_0_downstream_read;
  input            Medipix_sopc_burst_0_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_0_downstream_writedata;
  input   [ 10: 0] Medipix_sopc_burst_1_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_1_downstream_arbitrationshare;
  input            Medipix_sopc_burst_1_downstream_burstcount;
  input   [  3: 0] Medipix_sopc_burst_1_downstream_byteenable;
  input            Medipix_sopc_burst_1_downstream_debugaccess;
  input            Medipix_sopc_burst_1_downstream_latency_counter;
  input            Medipix_sopc_burst_1_downstream_read;
  input            Medipix_sopc_burst_1_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_1_downstream_writedata;
  input            clk;
  input   [ 31: 0] cpu_linux_jtag_debug_module_readdata;
  input            cpu_linux_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             Medipix_sopc_burst_0_downstream_arbiterlock;
  wire             Medipix_sopc_burst_0_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_0_downstream_continuerequest;
  wire             Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_saved_grant_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_arbiterlock;
  wire             Medipix_sopc_burst_1_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_1_downstream_continuerequest;
  wire             Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_saved_grant_cpu_linux_jtag_debug_module;
  wire    [  8: 0] cpu_linux_jtag_debug_module_address;
  wire             cpu_linux_jtag_debug_module_allgrants;
  wire             cpu_linux_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_linux_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_linux_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_linux_jtag_debug_module_arb_addend;
  wire             cpu_linux_jtag_debug_module_arb_counter_enable;
  reg     [  3: 0] cpu_linux_jtag_debug_module_arb_share_counter;
  wire    [  3: 0] cpu_linux_jtag_debug_module_arb_share_counter_next_value;
  wire    [  3: 0] cpu_linux_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_linux_jtag_debug_module_arb_winner;
  wire             cpu_linux_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_linux_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_linux_jtag_debug_module_begins_xfer;
  wire             cpu_linux_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_linux_jtag_debug_module_byteenable;
  wire             cpu_linux_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_linux_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_linux_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_linux_jtag_debug_module_debugaccess;
  wire             cpu_linux_jtag_debug_module_end_xfer;
  wire             cpu_linux_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_linux_jtag_debug_module_grant_vector;
  wire             cpu_linux_jtag_debug_module_in_a_read_cycle;
  wire             cpu_linux_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_linux_jtag_debug_module_master_qreq_vector;
  wire             cpu_linux_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_linux_jtag_debug_module_readdata_from_sa;
  reg              cpu_linux_jtag_debug_module_reg_firsttransfer;
  wire             cpu_linux_jtag_debug_module_reset_n;
  wire             cpu_linux_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_linux_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_linux_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_linux_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_linux_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_linux_jtag_debug_module_waits_for_read;
  wire             cpu_linux_jtag_debug_module_waits_for_write;
  wire             cpu_linux_jtag_debug_module_write;
  wire    [ 31: 0] cpu_linux_jtag_debug_module_writedata;
  reg              d1_cpu_linux_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_Medipix_sopc_burst_0_downstream_granted_slave_cpu_linux_jtag_debug_module;
  reg              last_cycle_Medipix_sopc_burst_1_downstream_granted_slave_cpu_linux_jtag_debug_module;
  wire    [ 10: 0] shifted_address_to_cpu_linux_jtag_debug_module_from_Medipix_sopc_burst_0_downstream;
  wire    [ 10: 0] shifted_address_to_cpu_linux_jtag_debug_module_from_Medipix_sopc_burst_1_downstream;
  wire             wait_for_cpu_linux_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_linux_jtag_debug_module_end_xfer;
    end


  assign cpu_linux_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module | Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module));
  //assign cpu_linux_jtag_debug_module_readdata_from_sa = cpu_linux_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_linux_jtag_debug_module_readdata_from_sa = cpu_linux_jtag_debug_module_readdata;

  assign Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module = (1) & (Medipix_sopc_burst_0_downstream_read | Medipix_sopc_burst_0_downstream_write);
  //cpu_linux_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_linux_jtag_debug_module_arb_share_set_values = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_0_downstream_arbitrationshare :
    (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_1_downstream_arbitrationshare :
    (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_0_downstream_arbitrationshare :
    (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_1_downstream_arbitrationshare :
    1;

  //cpu_linux_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_linux_jtag_debug_module_non_bursting_master_requests = 0;

  //cpu_linux_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_linux_jtag_debug_module_any_bursting_master_saved_grant = Medipix_sopc_burst_0_downstream_saved_grant_cpu_linux_jtag_debug_module |
    Medipix_sopc_burst_1_downstream_saved_grant_cpu_linux_jtag_debug_module |
    Medipix_sopc_burst_0_downstream_saved_grant_cpu_linux_jtag_debug_module |
    Medipix_sopc_burst_1_downstream_saved_grant_cpu_linux_jtag_debug_module;

  //cpu_linux_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_linux_jtag_debug_module_arb_share_counter_next_value = cpu_linux_jtag_debug_module_firsttransfer ? (cpu_linux_jtag_debug_module_arb_share_set_values - 1) : |cpu_linux_jtag_debug_module_arb_share_counter ? (cpu_linux_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_linux_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_linux_jtag_debug_module_allgrants = (|cpu_linux_jtag_debug_module_grant_vector) |
    (|cpu_linux_jtag_debug_module_grant_vector) |
    (|cpu_linux_jtag_debug_module_grant_vector) |
    (|cpu_linux_jtag_debug_module_grant_vector);

  //cpu_linux_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_linux_jtag_debug_module_end_xfer = ~(cpu_linux_jtag_debug_module_waits_for_read | cpu_linux_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module = cpu_linux_jtag_debug_module_end_xfer & (~cpu_linux_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_linux_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_linux_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module & cpu_linux_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module & ~cpu_linux_jtag_debug_module_non_bursting_master_requests);

  //cpu_linux_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_linux_jtag_debug_module_arb_counter_enable)
          cpu_linux_jtag_debug_module_arb_share_counter <= cpu_linux_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_linux_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_linux_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_linux_jtag_debug_module & ~cpu_linux_jtag_debug_module_non_bursting_master_requests))
          cpu_linux_jtag_debug_module_slavearbiterlockenable <= |cpu_linux_jtag_debug_module_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_0/downstream cpu_linux/jtag_debug_module arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_arbiterlock = cpu_linux_jtag_debug_module_slavearbiterlockenable & Medipix_sopc_burst_0_downstream_continuerequest;

  //cpu_linux_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_linux_jtag_debug_module_slavearbiterlockenable2 = |cpu_linux_jtag_debug_module_arb_share_counter_next_value;

  //Medipix_sopc_burst_0/downstream cpu_linux/jtag_debug_module arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_arbiterlock2 = cpu_linux_jtag_debug_module_slavearbiterlockenable2 & Medipix_sopc_burst_0_downstream_continuerequest;

  //Medipix_sopc_burst_1/downstream cpu_linux/jtag_debug_module arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_arbiterlock = cpu_linux_jtag_debug_module_slavearbiterlockenable & Medipix_sopc_burst_1_downstream_continuerequest;

  //Medipix_sopc_burst_1/downstream cpu_linux/jtag_debug_module arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_arbiterlock2 = cpu_linux_jtag_debug_module_slavearbiterlockenable2 & Medipix_sopc_burst_1_downstream_continuerequest;

  //Medipix_sopc_burst_1/downstream granted cpu_linux/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_Medipix_sopc_burst_1_downstream_granted_slave_cpu_linux_jtag_debug_module <= 0;
      else 
        last_cycle_Medipix_sopc_burst_1_downstream_granted_slave_cpu_linux_jtag_debug_module <= Medipix_sopc_burst_1_downstream_saved_grant_cpu_linux_jtag_debug_module ? 1 : (cpu_linux_jtag_debug_module_arbitration_holdoff_internal | 0) ? 0 : last_cycle_Medipix_sopc_burst_1_downstream_granted_slave_cpu_linux_jtag_debug_module;
    end


  //Medipix_sopc_burst_1_downstream_continuerequest continued request, which is an e_mux
  assign Medipix_sopc_burst_1_downstream_continuerequest = last_cycle_Medipix_sopc_burst_1_downstream_granted_slave_cpu_linux_jtag_debug_module & 1;

  //cpu_linux_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_linux_jtag_debug_module_any_continuerequest = Medipix_sopc_burst_1_downstream_continuerequest |
    Medipix_sopc_burst_0_downstream_continuerequest;

  assign Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module = Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module & ~((Medipix_sopc_burst_0_downstream_read & ((Medipix_sopc_burst_0_downstream_latency_counter != 0))) | Medipix_sopc_burst_1_downstream_arbiterlock);
  //local readdatavalid Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module, which is an e_mux
  assign Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module = Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_0_downstream_read & ~cpu_linux_jtag_debug_module_waits_for_read;

  //cpu_linux_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_linux_jtag_debug_module_writedata = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_0_downstream_writedata :
    Medipix_sopc_burst_1_downstream_writedata;

  assign Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module = (1) & (Medipix_sopc_burst_1_downstream_read | Medipix_sopc_burst_1_downstream_write);
  //Medipix_sopc_burst_0/downstream granted cpu_linux/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_Medipix_sopc_burst_0_downstream_granted_slave_cpu_linux_jtag_debug_module <= 0;
      else 
        last_cycle_Medipix_sopc_burst_0_downstream_granted_slave_cpu_linux_jtag_debug_module <= Medipix_sopc_burst_0_downstream_saved_grant_cpu_linux_jtag_debug_module ? 1 : (cpu_linux_jtag_debug_module_arbitration_holdoff_internal | 0) ? 0 : last_cycle_Medipix_sopc_burst_0_downstream_granted_slave_cpu_linux_jtag_debug_module;
    end


  //Medipix_sopc_burst_0_downstream_continuerequest continued request, which is an e_mux
  assign Medipix_sopc_burst_0_downstream_continuerequest = last_cycle_Medipix_sopc_burst_0_downstream_granted_slave_cpu_linux_jtag_debug_module & 1;

  assign Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module = Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module & ~((Medipix_sopc_burst_1_downstream_read & ((Medipix_sopc_burst_1_downstream_latency_counter != 0))) | Medipix_sopc_burst_0_downstream_arbiterlock);
  //local readdatavalid Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module, which is an e_mux
  assign Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module = Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_1_downstream_read & ~cpu_linux_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu_linux/jtag_debug_module, which is an e_assign
  assign cpu_linux_jtag_debug_module_allow_new_arb_cycle = ~Medipix_sopc_burst_0_downstream_arbiterlock & ~Medipix_sopc_burst_1_downstream_arbiterlock;

  //Medipix_sopc_burst_1/downstream assignment into master qualified-requests vector for cpu_linux/jtag_debug_module, which is an e_assign
  assign cpu_linux_jtag_debug_module_master_qreq_vector[0] = Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module;

  //Medipix_sopc_burst_1/downstream grant cpu_linux/jtag_debug_module, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module = cpu_linux_jtag_debug_module_grant_vector[0];

  //Medipix_sopc_burst_1/downstream saved-grant cpu_linux/jtag_debug_module, which is an e_assign
  assign Medipix_sopc_burst_1_downstream_saved_grant_cpu_linux_jtag_debug_module = cpu_linux_jtag_debug_module_arb_winner[0];

  //Medipix_sopc_burst_0/downstream assignment into master qualified-requests vector for cpu_linux/jtag_debug_module, which is an e_assign
  assign cpu_linux_jtag_debug_module_master_qreq_vector[1] = Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module;

  //Medipix_sopc_burst_0/downstream grant cpu_linux/jtag_debug_module, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module = cpu_linux_jtag_debug_module_grant_vector[1];

  //Medipix_sopc_burst_0/downstream saved-grant cpu_linux/jtag_debug_module, which is an e_assign
  assign Medipix_sopc_burst_0_downstream_saved_grant_cpu_linux_jtag_debug_module = cpu_linux_jtag_debug_module_arb_winner[1];

  //cpu_linux/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_linux_jtag_debug_module_chosen_master_double_vector = {cpu_linux_jtag_debug_module_master_qreq_vector, cpu_linux_jtag_debug_module_master_qreq_vector} & ({~cpu_linux_jtag_debug_module_master_qreq_vector, ~cpu_linux_jtag_debug_module_master_qreq_vector} + cpu_linux_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_linux_jtag_debug_module_arb_winner = (cpu_linux_jtag_debug_module_allow_new_arb_cycle & | cpu_linux_jtag_debug_module_grant_vector) ? cpu_linux_jtag_debug_module_grant_vector : cpu_linux_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_linux_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_linux_jtag_debug_module_allow_new_arb_cycle)
          cpu_linux_jtag_debug_module_saved_chosen_master_vector <= |cpu_linux_jtag_debug_module_grant_vector ? cpu_linux_jtag_debug_module_grant_vector : cpu_linux_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_linux_jtag_debug_module_grant_vector = {(cpu_linux_jtag_debug_module_chosen_master_double_vector[1] | cpu_linux_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_linux_jtag_debug_module_chosen_master_double_vector[0] | cpu_linux_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu_linux/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_linux_jtag_debug_module_chosen_master_rot_left = (cpu_linux_jtag_debug_module_arb_winner << 1) ? (cpu_linux_jtag_debug_module_arb_winner << 1) : 1;

  //cpu_linux/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_linux_jtag_debug_module_grant_vector)
          cpu_linux_jtag_debug_module_arb_addend <= cpu_linux_jtag_debug_module_end_xfer? cpu_linux_jtag_debug_module_chosen_master_rot_left : cpu_linux_jtag_debug_module_grant_vector;
    end


  assign cpu_linux_jtag_debug_module_begintransfer = cpu_linux_jtag_debug_module_begins_xfer;
  //cpu_linux_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_linux_jtag_debug_module_reset_n = reset_n;

  //assign cpu_linux_jtag_debug_module_resetrequest_from_sa = cpu_linux_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_linux_jtag_debug_module_resetrequest_from_sa = cpu_linux_jtag_debug_module_resetrequest;

  assign cpu_linux_jtag_debug_module_chipselect = Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module | Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module;
  //cpu_linux_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_linux_jtag_debug_module_firsttransfer = cpu_linux_jtag_debug_module_begins_xfer ? cpu_linux_jtag_debug_module_unreg_firsttransfer : cpu_linux_jtag_debug_module_reg_firsttransfer;

  //cpu_linux_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_linux_jtag_debug_module_unreg_firsttransfer = ~(cpu_linux_jtag_debug_module_slavearbiterlockenable & cpu_linux_jtag_debug_module_any_continuerequest);

  //cpu_linux_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_linux_jtag_debug_module_begins_xfer)
          cpu_linux_jtag_debug_module_reg_firsttransfer <= cpu_linux_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_linux_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_linux_jtag_debug_module_beginbursttransfer_internal = cpu_linux_jtag_debug_module_begins_xfer;

  //cpu_linux_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_linux_jtag_debug_module_arbitration_holdoff_internal = cpu_linux_jtag_debug_module_begins_xfer & cpu_linux_jtag_debug_module_firsttransfer;

  //cpu_linux_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_linux_jtag_debug_module_write = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_0_downstream_write) | (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_1_downstream_write);

  assign shifted_address_to_cpu_linux_jtag_debug_module_from_Medipix_sopc_burst_0_downstream = Medipix_sopc_burst_0_downstream_address_to_slave;
  //cpu_linux_jtag_debug_module_address mux, which is an e_mux
  assign cpu_linux_jtag_debug_module_address = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module)? (shifted_address_to_cpu_linux_jtag_debug_module_from_Medipix_sopc_burst_0_downstream >> 2) :
    (shifted_address_to_cpu_linux_jtag_debug_module_from_Medipix_sopc_burst_1_downstream >> 2);

  assign shifted_address_to_cpu_linux_jtag_debug_module_from_Medipix_sopc_burst_1_downstream = Medipix_sopc_burst_1_downstream_address_to_slave;
  //d1_cpu_linux_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_linux_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_linux_jtag_debug_module_end_xfer <= cpu_linux_jtag_debug_module_end_xfer;
    end


  //cpu_linux_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_linux_jtag_debug_module_waits_for_read = cpu_linux_jtag_debug_module_in_a_read_cycle & cpu_linux_jtag_debug_module_begins_xfer;

  //cpu_linux_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_linux_jtag_debug_module_in_a_read_cycle = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_0_downstream_read) | (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_1_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_linux_jtag_debug_module_in_a_read_cycle;

  //cpu_linux_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_linux_jtag_debug_module_waits_for_write = cpu_linux_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_linux_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_linux_jtag_debug_module_in_a_write_cycle = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_0_downstream_write) | (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module & Medipix_sopc_burst_1_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_linux_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_linux_jtag_debug_module_counter = 0;
  //cpu_linux_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_linux_jtag_debug_module_byteenable = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_0_downstream_byteenable :
    (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_1_downstream_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_linux_jtag_debug_module_debugaccess = (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_0_downstream_debugaccess :
    (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module)? Medipix_sopc_burst_1_downstream_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_linux/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module && (Medipix_sopc_burst_0_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave cpu_linux/jtag_debug_module", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_0/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module && (Medipix_sopc_burst_0_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave cpu_linux/jtag_debug_module", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module && (Medipix_sopc_burst_1_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_1/downstream drove 0 on its 'arbitrationshare' port while accessing slave cpu_linux/jtag_debug_module", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_1/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module && (Medipix_sopc_burst_1_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_1/downstream drove 0 on its 'burstcount' port while accessing slave cpu_linux/jtag_debug_module", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module + Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_0_downstream_saved_grant_cpu_linux_jtag_debug_module + Medipix_sopc_burst_1_downstream_saved_grant_cpu_linux_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_linux_data_master_arbitrator (
                                          // inputs:
                                           Medipix_sopc_burst_10_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_10_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_11_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_11_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_1_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_1_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_2_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_2_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_3_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_3_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_5_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_5_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_7_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_7_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_8_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_8_upstream_waitrequest_from_sa,
                                           Medipix_sopc_burst_9_upstream_readdata_from_sa,
                                           Medipix_sopc_burst_9_upstream_waitrequest_from_sa,
                                           clk,
                                           cpu_linux_data_master_address,
                                           cpu_linux_data_master_burstcount,
                                           cpu_linux_data_master_byteenable,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream,
                                           cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream,
                                           cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream,
                                           cpu_linux_data_master_read,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream,
                                           cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream,
                                           cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream,
                                           cpu_linux_data_master_write,
                                           cpu_linux_data_master_writedata,
                                           d1_Medipix_sopc_burst_10_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_11_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_1_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_2_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_3_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_5_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_7_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_8_upstream_end_xfer,
                                           d1_Medipix_sopc_burst_9_upstream_end_xfer,
                                           epcs_controller_epcs_control_port_irq_from_sa,
                                           igor_mac_control_port_irq_from_sa,
                                           jtag_uart_0_avalon_jtag_slave_irq_from_sa,
                                           reset_n,
                                           spi_0_spi_control_port_irq_from_sa,
                                           sys_clk_freq_s1_irq_from_sa,
                                           uart_0_s1_irq_from_sa,

                                          // outputs:
                                           cpu_linux_data_master_address_to_slave,
                                           cpu_linux_data_master_irq,
                                           cpu_linux_data_master_latency_counter,
                                           cpu_linux_data_master_readdata,
                                           cpu_linux_data_master_readdatavalid,
                                           cpu_linux_data_master_waitrequest
                                        )
;

  output  [ 27: 0] cpu_linux_data_master_address_to_slave;
  output  [ 31: 0] cpu_linux_data_master_irq;
  output           cpu_linux_data_master_latency_counter;
  output  [ 31: 0] cpu_linux_data_master_readdata;
  output           cpu_linux_data_master_readdatavalid;
  output           cpu_linux_data_master_waitrequest;
  input   [ 15: 0] Medipix_sopc_burst_10_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_10_upstream_waitrequest_from_sa;
  input   [ 15: 0] Medipix_sopc_burst_11_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_11_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_1_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_1_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_2_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_2_upstream_waitrequest_from_sa;
  input   [ 15: 0] Medipix_sopc_burst_3_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_3_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_5_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_5_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_7_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_7_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_8_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_8_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_9_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_9_upstream_waitrequest_from_sa;
  input            clk;
  input   [ 27: 0] cpu_linux_data_master_address;
  input   [  3: 0] cpu_linux_data_master_burstcount;
  input   [  3: 0] cpu_linux_data_master_byteenable;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream;
  input            cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream;
  input            cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream;
  input            cpu_linux_data_master_read;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream;
  input            cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream;
  input            cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream;
  input            cpu_linux_data_master_write;
  input   [ 31: 0] cpu_linux_data_master_writedata;
  input            d1_Medipix_sopc_burst_10_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_11_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_1_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_2_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_3_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_5_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_7_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_8_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_9_upstream_end_xfer;
  input            epcs_controller_epcs_control_port_irq_from_sa;
  input            igor_mac_control_port_irq_from_sa;
  input            jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  input            reset_n;
  input            spi_0_spi_control_port_irq_from_sa;
  input            sys_clk_freq_s1_irq_from_sa;
  input            uart_0_s1_irq_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 27: 0] cpu_linux_data_master_address_last_time;
  wire    [ 27: 0] cpu_linux_data_master_address_to_slave;
  reg     [  3: 0] cpu_linux_data_master_burstcount_last_time;
  reg     [  3: 0] cpu_linux_data_master_byteenable_last_time;
  wire    [ 31: 0] cpu_linux_data_master_irq;
  wire             cpu_linux_data_master_is_granted_some_slave;
  reg              cpu_linux_data_master_latency_counter;
  reg              cpu_linux_data_master_read_but_no_slave_selected;
  reg              cpu_linux_data_master_read_last_time;
  wire    [ 31: 0] cpu_linux_data_master_readdata;
  wire             cpu_linux_data_master_readdatavalid;
  wire             cpu_linux_data_master_run;
  wire             cpu_linux_data_master_waitrequest;
  reg              cpu_linux_data_master_write_last_time;
  reg     [ 31: 0] cpu_linux_data_master_writedata_last_time;
  wire             latency_load_value;
  wire             p1_cpu_linux_data_master_latency_counter;
  wire             pre_flush_cpu_linux_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_1_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_1_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_10_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_10_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_11_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_11_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_2_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_2_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_3_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_3_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_linux_data_master_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_5_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_5_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_7_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_7_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_8_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_8_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & 1 & (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream | ~cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_9_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write)))) & ((~cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream | ~(cpu_linux_data_master_read | cpu_linux_data_master_write) | (1 & ~Medipix_sopc_burst_9_upstream_waitrequest_from_sa & (cpu_linux_data_master_read | cpu_linux_data_master_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_linux_data_master_address_to_slave = cpu_linux_data_master_address[27 : 0];

  //cpu_linux_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_linux_data_master_read_but_no_slave_selected <= cpu_linux_data_master_read & cpu_linux_data_master_run & ~cpu_linux_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_linux_data_master_is_granted_some_slave = cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream |
    cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_linux_data_master_readdatavalid = cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream |
    cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_linux_data_master_readdatavalid = cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid |
    cpu_linux_data_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_data_master_readdatavalid;

  //cpu_linux/data_master readdata mux, which is an e_mux
  assign cpu_linux_data_master_readdata = ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream}} | Medipix_sopc_burst_1_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream}} | Medipix_sopc_burst_10_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream}} | Medipix_sopc_burst_11_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream}} | Medipix_sopc_burst_2_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream}} | Medipix_sopc_burst_3_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream}} | Medipix_sopc_burst_5_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream}} | Medipix_sopc_burst_7_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream}} | Medipix_sopc_burst_8_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream}} | Medipix_sopc_burst_9_upstream_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_linux_data_master_waitrequest = ~cpu_linux_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_latency_counter <= 0;
      else 
        cpu_linux_data_master_latency_counter <= p1_cpu_linux_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_linux_data_master_latency_counter = ((cpu_linux_data_master_run & cpu_linux_data_master_read))? latency_load_value :
    (cpu_linux_data_master_latency_counter)? cpu_linux_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //irq assign, which is an e_assign
  assign cpu_linux_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    spi_0_spi_control_port_irq_from_sa,
    uart_0_s1_irq_from_sa,
    igor_mac_control_port_irq_from_sa,
    epcs_controller_epcs_control_port_irq_from_sa,
    jtag_uart_0_avalon_jtag_slave_irq_from_sa,
    sys_clk_freq_s1_irq_from_sa};


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_linux_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_address_last_time <= 0;
      else 
        cpu_linux_data_master_address_last_time <= cpu_linux_data_master_address;
    end


  //cpu_linux/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_linux_data_master_waitrequest & (cpu_linux_data_master_read | cpu_linux_data_master_write);
    end


  //cpu_linux_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_data_master_address != cpu_linux_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_linux_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_data_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_burstcount_last_time <= 0;
      else 
        cpu_linux_data_master_burstcount_last_time <= cpu_linux_data_master_burstcount;
    end


  //cpu_linux_data_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_data_master_burstcount != cpu_linux_data_master_burstcount_last_time))
        begin
          $write("%0d ns: cpu_linux_data_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_byteenable_last_time <= 0;
      else 
        cpu_linux_data_master_byteenable_last_time <= cpu_linux_data_master_byteenable;
    end


  //cpu_linux_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_data_master_byteenable != cpu_linux_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_linux_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_read_last_time <= 0;
      else 
        cpu_linux_data_master_read_last_time <= cpu_linux_data_master_read;
    end


  //cpu_linux_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_data_master_read != cpu_linux_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_linux_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_write_last_time <= 0;
      else 
        cpu_linux_data_master_write_last_time <= cpu_linux_data_master_write;
    end


  //cpu_linux_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_data_master_write != cpu_linux_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_linux_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_data_master_writedata_last_time <= 0;
      else 
        cpu_linux_data_master_writedata_last_time <= cpu_linux_data_master_writedata;
    end


  //cpu_linux_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_data_master_writedata != cpu_linux_data_master_writedata_last_time) & cpu_linux_data_master_write)
        begin
          $write("%0d ns: cpu_linux_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_linux_instruction_master_arbitrator (
                                                 // inputs:
                                                  Medipix_sopc_burst_0_upstream_readdata_from_sa,
                                                  Medipix_sopc_burst_0_upstream_waitrequest_from_sa,
                                                  Medipix_sopc_burst_4_upstream_readdata_from_sa,
                                                  Medipix_sopc_burst_4_upstream_waitrequest_from_sa,
                                                  Medipix_sopc_burst_6_upstream_readdata_from_sa,
                                                  Medipix_sopc_burst_6_upstream_waitrequest_from_sa,
                                                  clk,
                                                  cpu_linux_instruction_master_address,
                                                  cpu_linux_instruction_master_burstcount,
                                                  cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream,
                                                  cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream,
                                                  cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream,
                                                  cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream,
                                                  cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream,
                                                  cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream,
                                                  cpu_linux_instruction_master_read,
                                                  cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream,
                                                  cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register,
                                                  cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream,
                                                  cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register,
                                                  cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream,
                                                  cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register,
                                                  cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream,
                                                  cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream,
                                                  cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream,
                                                  d1_Medipix_sopc_burst_0_upstream_end_xfer,
                                                  d1_Medipix_sopc_burst_4_upstream_end_xfer,
                                                  d1_Medipix_sopc_burst_6_upstream_end_xfer,
                                                  reset_n,

                                                 // outputs:
                                                  cpu_linux_instruction_master_address_to_slave,
                                                  cpu_linux_instruction_master_latency_counter,
                                                  cpu_linux_instruction_master_readdata,
                                                  cpu_linux_instruction_master_readdatavalid,
                                                  cpu_linux_instruction_master_waitrequest
                                               )
;

  output  [ 27: 0] cpu_linux_instruction_master_address_to_slave;
  output           cpu_linux_instruction_master_latency_counter;
  output  [ 31: 0] cpu_linux_instruction_master_readdata;
  output           cpu_linux_instruction_master_readdatavalid;
  output           cpu_linux_instruction_master_waitrequest;
  input   [ 31: 0] Medipix_sopc_burst_0_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_0_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_4_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_4_upstream_waitrequest_from_sa;
  input   [ 31: 0] Medipix_sopc_burst_6_upstream_readdata_from_sa;
  input            Medipix_sopc_burst_6_upstream_waitrequest_from_sa;
  input            clk;
  input   [ 27: 0] cpu_linux_instruction_master_address;
  input   [  3: 0] cpu_linux_instruction_master_burstcount;
  input            cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream;
  input            cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream;
  input            cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream;
  input            cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream;
  input            cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream;
  input            cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream;
  input            cpu_linux_instruction_master_read;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream;
  input            cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register;
  input            cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream;
  input            cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream;
  input            cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream;
  input            d1_Medipix_sopc_burst_0_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_4_upstream_end_xfer;
  input            d1_Medipix_sopc_burst_6_upstream_end_xfer;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 27: 0] cpu_linux_instruction_master_address_last_time;
  wire    [ 27: 0] cpu_linux_instruction_master_address_to_slave;
  reg     [  3: 0] cpu_linux_instruction_master_burstcount_last_time;
  wire             cpu_linux_instruction_master_is_granted_some_slave;
  reg              cpu_linux_instruction_master_latency_counter;
  reg              cpu_linux_instruction_master_read_but_no_slave_selected;
  reg              cpu_linux_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_linux_instruction_master_readdata;
  wire             cpu_linux_instruction_master_readdatavalid;
  wire             cpu_linux_instruction_master_run;
  wire             cpu_linux_instruction_master_waitrequest;
  wire             latency_load_value;
  wire             p1_cpu_linux_instruction_master_latency_counter;
  wire             pre_flush_cpu_linux_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream | ~cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream) & ((~cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream | ~(cpu_linux_instruction_master_read) | (1 & ~Medipix_sopc_burst_0_upstream_waitrequest_from_sa & (cpu_linux_instruction_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_linux_instruction_master_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream | ~cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream) & ((~cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream | ~(cpu_linux_instruction_master_read) | (1 & ~Medipix_sopc_burst_4_upstream_waitrequest_from_sa & (cpu_linux_instruction_master_read)))) & 1 & (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream | ~cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream) & ((~cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream | ~(cpu_linux_instruction_master_read) | (1 & ~Medipix_sopc_burst_6_upstream_waitrequest_from_sa & (cpu_linux_instruction_master_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_linux_instruction_master_address_to_slave = cpu_linux_instruction_master_address[27 : 0];

  //cpu_linux_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_linux_instruction_master_read_but_no_slave_selected <= cpu_linux_instruction_master_read & cpu_linux_instruction_master_run & ~cpu_linux_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_linux_instruction_master_is_granted_some_slave = cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream |
    cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream |
    cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_linux_instruction_master_readdatavalid = cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream |
    cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream |
    cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_linux_instruction_master_readdatavalid = cpu_linux_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_instruction_master_readdatavalid |
    cpu_linux_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_instruction_master_readdatavalid |
    cpu_linux_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_linux_instruction_master_readdatavalid;

  //cpu_linux/instruction_master readdata mux, which is an e_mux
  assign cpu_linux_instruction_master_readdata = ({32 {~cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream}} | Medipix_sopc_burst_0_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream}} | Medipix_sopc_burst_4_upstream_readdata_from_sa) &
    ({32 {~cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream}} | Medipix_sopc_burst_6_upstream_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_linux_instruction_master_waitrequest = ~cpu_linux_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_instruction_master_latency_counter <= 0;
      else 
        cpu_linux_instruction_master_latency_counter <= p1_cpu_linux_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_linux_instruction_master_latency_counter = ((cpu_linux_instruction_master_run & cpu_linux_instruction_master_read))? latency_load_value :
    (cpu_linux_instruction_master_latency_counter)? cpu_linux_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_linux_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_instruction_master_address_last_time <= 0;
      else 
        cpu_linux_instruction_master_address_last_time <= cpu_linux_instruction_master_address;
    end


  //cpu_linux/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_linux_instruction_master_waitrequest & (cpu_linux_instruction_master_read);
    end


  //cpu_linux_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_instruction_master_address != cpu_linux_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_linux_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_instruction_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_instruction_master_burstcount_last_time <= 0;
      else 
        cpu_linux_instruction_master_burstcount_last_time <= cpu_linux_instruction_master_burstcount;
    end


  //cpu_linux_instruction_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_instruction_master_burstcount != cpu_linux_instruction_master_burstcount_last_time))
        begin
          $write("%0d ns: cpu_linux_instruction_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_linux_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_linux_instruction_master_read_last_time <= 0;
      else 
        cpu_linux_instruction_master_read_last_time <= cpu_linux_instruction_master_read;
    end


  //cpu_linux_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_linux_instruction_master_read != cpu_linux_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_linux_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module epcs_controller_epcs_control_port_arbitrator (
                                                      // inputs:
                                                       Medipix_sopc_burst_6_downstream_address_to_slave,
                                                       Medipix_sopc_burst_6_downstream_arbitrationshare,
                                                       Medipix_sopc_burst_6_downstream_burstcount,
                                                       Medipix_sopc_burst_6_downstream_latency_counter,
                                                       Medipix_sopc_burst_6_downstream_read,
                                                       Medipix_sopc_burst_6_downstream_write,
                                                       Medipix_sopc_burst_6_downstream_writedata,
                                                       Medipix_sopc_burst_7_downstream_address_to_slave,
                                                       Medipix_sopc_burst_7_downstream_arbitrationshare,
                                                       Medipix_sopc_burst_7_downstream_burstcount,
                                                       Medipix_sopc_burst_7_downstream_latency_counter,
                                                       Medipix_sopc_burst_7_downstream_read,
                                                       Medipix_sopc_burst_7_downstream_write,
                                                       Medipix_sopc_burst_7_downstream_writedata,
                                                       clk,
                                                       epcs_controller_epcs_control_port_dataavailable,
                                                       epcs_controller_epcs_control_port_endofpacket,
                                                       epcs_controller_epcs_control_port_irq,
                                                       epcs_controller_epcs_control_port_readdata,
                                                       epcs_controller_epcs_control_port_readyfordata,
                                                       reset_n,

                                                      // outputs:
                                                       Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port,
                                                       Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port,
                                                       d1_epcs_controller_epcs_control_port_end_xfer,
                                                       epcs_controller_epcs_control_port_address,
                                                       epcs_controller_epcs_control_port_chipselect,
                                                       epcs_controller_epcs_control_port_dataavailable_from_sa,
                                                       epcs_controller_epcs_control_port_endofpacket_from_sa,
                                                       epcs_controller_epcs_control_port_irq_from_sa,
                                                       epcs_controller_epcs_control_port_read_n,
                                                       epcs_controller_epcs_control_port_readdata_from_sa,
                                                       epcs_controller_epcs_control_port_readyfordata_from_sa,
                                                       epcs_controller_epcs_control_port_reset_n,
                                                       epcs_controller_epcs_control_port_write_n,
                                                       epcs_controller_epcs_control_port_writedata
                                                    )
;

  output           Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port;
  output           Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port;
  output           d1_epcs_controller_epcs_control_port_end_xfer;
  output  [  8: 0] epcs_controller_epcs_control_port_address;
  output           epcs_controller_epcs_control_port_chipselect;
  output           epcs_controller_epcs_control_port_dataavailable_from_sa;
  output           epcs_controller_epcs_control_port_endofpacket_from_sa;
  output           epcs_controller_epcs_control_port_irq_from_sa;
  output           epcs_controller_epcs_control_port_read_n;
  output  [ 31: 0] epcs_controller_epcs_control_port_readdata_from_sa;
  output           epcs_controller_epcs_control_port_readyfordata_from_sa;
  output           epcs_controller_epcs_control_port_reset_n;
  output           epcs_controller_epcs_control_port_write_n;
  output  [ 31: 0] epcs_controller_epcs_control_port_writedata;
  input   [ 10: 0] Medipix_sopc_burst_6_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_6_downstream_arbitrationshare;
  input            Medipix_sopc_burst_6_downstream_burstcount;
  input            Medipix_sopc_burst_6_downstream_latency_counter;
  input            Medipix_sopc_burst_6_downstream_read;
  input            Medipix_sopc_burst_6_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_6_downstream_writedata;
  input   [ 10: 0] Medipix_sopc_burst_7_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_7_downstream_arbitrationshare;
  input            Medipix_sopc_burst_7_downstream_burstcount;
  input            Medipix_sopc_burst_7_downstream_latency_counter;
  input            Medipix_sopc_burst_7_downstream_read;
  input            Medipix_sopc_burst_7_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_7_downstream_writedata;
  input            clk;
  input            epcs_controller_epcs_control_port_dataavailable;
  input            epcs_controller_epcs_control_port_endofpacket;
  input            epcs_controller_epcs_control_port_irq;
  input   [ 31: 0] epcs_controller_epcs_control_port_readdata;
  input            epcs_controller_epcs_control_port_readyfordata;
  input            reset_n;

  wire             Medipix_sopc_burst_6_downstream_arbiterlock;
  wire             Medipix_sopc_burst_6_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_6_downstream_continuerequest;
  wire             Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_saved_grant_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_arbiterlock;
  wire             Medipix_sopc_burst_7_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_7_downstream_continuerequest;
  wire             Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_saved_grant_epcs_controller_epcs_control_port;
  reg              d1_epcs_controller_epcs_control_port_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port;
  wire    [  8: 0] epcs_controller_epcs_control_port_address;
  wire             epcs_controller_epcs_control_port_allgrants;
  wire             epcs_controller_epcs_control_port_allow_new_arb_cycle;
  wire             epcs_controller_epcs_control_port_any_bursting_master_saved_grant;
  wire             epcs_controller_epcs_control_port_any_continuerequest;
  reg     [  1: 0] epcs_controller_epcs_control_port_arb_addend;
  wire             epcs_controller_epcs_control_port_arb_counter_enable;
  reg     [  3: 0] epcs_controller_epcs_control_port_arb_share_counter;
  wire    [  3: 0] epcs_controller_epcs_control_port_arb_share_counter_next_value;
  wire    [  3: 0] epcs_controller_epcs_control_port_arb_share_set_values;
  wire    [  1: 0] epcs_controller_epcs_control_port_arb_winner;
  wire             epcs_controller_epcs_control_port_arbitration_holdoff_internal;
  wire             epcs_controller_epcs_control_port_beginbursttransfer_internal;
  wire             epcs_controller_epcs_control_port_begins_xfer;
  wire             epcs_controller_epcs_control_port_chipselect;
  wire    [  3: 0] epcs_controller_epcs_control_port_chosen_master_double_vector;
  wire    [  1: 0] epcs_controller_epcs_control_port_chosen_master_rot_left;
  wire             epcs_controller_epcs_control_port_dataavailable_from_sa;
  wire             epcs_controller_epcs_control_port_end_xfer;
  wire             epcs_controller_epcs_control_port_endofpacket_from_sa;
  wire             epcs_controller_epcs_control_port_firsttransfer;
  wire    [  1: 0] epcs_controller_epcs_control_port_grant_vector;
  wire             epcs_controller_epcs_control_port_in_a_read_cycle;
  wire             epcs_controller_epcs_control_port_in_a_write_cycle;
  wire             epcs_controller_epcs_control_port_irq_from_sa;
  wire    [  1: 0] epcs_controller_epcs_control_port_master_qreq_vector;
  wire             epcs_controller_epcs_control_port_non_bursting_master_requests;
  wire             epcs_controller_epcs_control_port_read_n;
  wire    [ 31: 0] epcs_controller_epcs_control_port_readdata_from_sa;
  wire             epcs_controller_epcs_control_port_readyfordata_from_sa;
  reg              epcs_controller_epcs_control_port_reg_firsttransfer;
  wire             epcs_controller_epcs_control_port_reset_n;
  reg     [  1: 0] epcs_controller_epcs_control_port_saved_chosen_master_vector;
  reg              epcs_controller_epcs_control_port_slavearbiterlockenable;
  wire             epcs_controller_epcs_control_port_slavearbiterlockenable2;
  wire             epcs_controller_epcs_control_port_unreg_firsttransfer;
  wire             epcs_controller_epcs_control_port_waits_for_read;
  wire             epcs_controller_epcs_control_port_waits_for_write;
  wire             epcs_controller_epcs_control_port_write_n;
  wire    [ 31: 0] epcs_controller_epcs_control_port_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_Medipix_sopc_burst_6_downstream_granted_slave_epcs_controller_epcs_control_port;
  reg              last_cycle_Medipix_sopc_burst_7_downstream_granted_slave_epcs_controller_epcs_control_port;
  wire    [ 10: 0] shifted_address_to_epcs_controller_epcs_control_port_from_Medipix_sopc_burst_6_downstream;
  wire    [ 10: 0] shifted_address_to_epcs_controller_epcs_control_port_from_Medipix_sopc_burst_7_downstream;
  wire             wait_for_epcs_controller_epcs_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~epcs_controller_epcs_control_port_end_xfer;
    end


  assign epcs_controller_epcs_control_port_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port | Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port));
  //assign epcs_controller_epcs_control_port_readdata_from_sa = epcs_controller_epcs_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_controller_epcs_control_port_readdata_from_sa = epcs_controller_epcs_control_port_readdata;

  assign Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port = (1) & (Medipix_sopc_burst_6_downstream_read | Medipix_sopc_burst_6_downstream_write);
  //assign epcs_controller_epcs_control_port_dataavailable_from_sa = epcs_controller_epcs_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_controller_epcs_control_port_dataavailable_from_sa = epcs_controller_epcs_control_port_dataavailable;

  //assign epcs_controller_epcs_control_port_readyfordata_from_sa = epcs_controller_epcs_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_controller_epcs_control_port_readyfordata_from_sa = epcs_controller_epcs_control_port_readyfordata;

  //epcs_controller_epcs_control_port_arb_share_counter set values, which is an e_mux
  assign epcs_controller_epcs_control_port_arb_share_set_values = (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port)? Medipix_sopc_burst_6_downstream_arbitrationshare :
    (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port)? Medipix_sopc_burst_7_downstream_arbitrationshare :
    (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port)? Medipix_sopc_burst_6_downstream_arbitrationshare :
    (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port)? Medipix_sopc_burst_7_downstream_arbitrationshare :
    1;

  //epcs_controller_epcs_control_port_non_bursting_master_requests mux, which is an e_mux
  assign epcs_controller_epcs_control_port_non_bursting_master_requests = 0;

  //epcs_controller_epcs_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign epcs_controller_epcs_control_port_any_bursting_master_saved_grant = Medipix_sopc_burst_6_downstream_saved_grant_epcs_controller_epcs_control_port |
    Medipix_sopc_burst_7_downstream_saved_grant_epcs_controller_epcs_control_port |
    Medipix_sopc_burst_6_downstream_saved_grant_epcs_controller_epcs_control_port |
    Medipix_sopc_burst_7_downstream_saved_grant_epcs_controller_epcs_control_port;

  //epcs_controller_epcs_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign epcs_controller_epcs_control_port_arb_share_counter_next_value = epcs_controller_epcs_control_port_firsttransfer ? (epcs_controller_epcs_control_port_arb_share_set_values - 1) : |epcs_controller_epcs_control_port_arb_share_counter ? (epcs_controller_epcs_control_port_arb_share_counter - 1) : 0;

  //epcs_controller_epcs_control_port_allgrants all slave grants, which is an e_mux
  assign epcs_controller_epcs_control_port_allgrants = (|epcs_controller_epcs_control_port_grant_vector) |
    (|epcs_controller_epcs_control_port_grant_vector) |
    (|epcs_controller_epcs_control_port_grant_vector) |
    (|epcs_controller_epcs_control_port_grant_vector);

  //epcs_controller_epcs_control_port_end_xfer assignment, which is an e_assign
  assign epcs_controller_epcs_control_port_end_xfer = ~(epcs_controller_epcs_control_port_waits_for_read | epcs_controller_epcs_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port = epcs_controller_epcs_control_port_end_xfer & (~epcs_controller_epcs_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //epcs_controller_epcs_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign epcs_controller_epcs_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port & epcs_controller_epcs_control_port_allgrants) | (end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port & ~epcs_controller_epcs_control_port_non_bursting_master_requests);

  //epcs_controller_epcs_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_controller_epcs_control_port_arb_share_counter <= 0;
      else if (epcs_controller_epcs_control_port_arb_counter_enable)
          epcs_controller_epcs_control_port_arb_share_counter <= epcs_controller_epcs_control_port_arb_share_counter_next_value;
    end


  //epcs_controller_epcs_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_controller_epcs_control_port_slavearbiterlockenable <= 0;
      else if ((|epcs_controller_epcs_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port) | (end_xfer_arb_share_counter_term_epcs_controller_epcs_control_port & ~epcs_controller_epcs_control_port_non_bursting_master_requests))
          epcs_controller_epcs_control_port_slavearbiterlockenable <= |epcs_controller_epcs_control_port_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_6/downstream epcs_controller/epcs_control_port arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_arbiterlock = epcs_controller_epcs_control_port_slavearbiterlockenable & Medipix_sopc_burst_6_downstream_continuerequest;

  //epcs_controller_epcs_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign epcs_controller_epcs_control_port_slavearbiterlockenable2 = |epcs_controller_epcs_control_port_arb_share_counter_next_value;

  //Medipix_sopc_burst_6/downstream epcs_controller/epcs_control_port arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_arbiterlock2 = epcs_controller_epcs_control_port_slavearbiterlockenable2 & Medipix_sopc_burst_6_downstream_continuerequest;

  //Medipix_sopc_burst_7/downstream epcs_controller/epcs_control_port arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_arbiterlock = epcs_controller_epcs_control_port_slavearbiterlockenable & Medipix_sopc_burst_7_downstream_continuerequest;

  //Medipix_sopc_burst_7/downstream epcs_controller/epcs_control_port arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_arbiterlock2 = epcs_controller_epcs_control_port_slavearbiterlockenable2 & Medipix_sopc_burst_7_downstream_continuerequest;

  //Medipix_sopc_burst_7/downstream granted epcs_controller/epcs_control_port last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_Medipix_sopc_burst_7_downstream_granted_slave_epcs_controller_epcs_control_port <= 0;
      else 
        last_cycle_Medipix_sopc_burst_7_downstream_granted_slave_epcs_controller_epcs_control_port <= Medipix_sopc_burst_7_downstream_saved_grant_epcs_controller_epcs_control_port ? 1 : (epcs_controller_epcs_control_port_arbitration_holdoff_internal | 0) ? 0 : last_cycle_Medipix_sopc_burst_7_downstream_granted_slave_epcs_controller_epcs_control_port;
    end


  //Medipix_sopc_burst_7_downstream_continuerequest continued request, which is an e_mux
  assign Medipix_sopc_burst_7_downstream_continuerequest = last_cycle_Medipix_sopc_burst_7_downstream_granted_slave_epcs_controller_epcs_control_port & 1;

  //epcs_controller_epcs_control_port_any_continuerequest at least one master continues requesting, which is an e_mux
  assign epcs_controller_epcs_control_port_any_continuerequest = Medipix_sopc_burst_7_downstream_continuerequest |
    Medipix_sopc_burst_6_downstream_continuerequest;

  assign Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port = Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port & ~((Medipix_sopc_burst_6_downstream_read & ((Medipix_sopc_burst_6_downstream_latency_counter != 0))) | Medipix_sopc_burst_7_downstream_arbiterlock);
  //local readdatavalid Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port, which is an e_mux
  assign Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port = Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_6_downstream_read & ~epcs_controller_epcs_control_port_waits_for_read;

  //epcs_controller_epcs_control_port_writedata mux, which is an e_mux
  assign epcs_controller_epcs_control_port_writedata = (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port)? Medipix_sopc_burst_6_downstream_writedata :
    Medipix_sopc_burst_7_downstream_writedata;

  //assign epcs_controller_epcs_control_port_endofpacket_from_sa = epcs_controller_epcs_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_controller_epcs_control_port_endofpacket_from_sa = epcs_controller_epcs_control_port_endofpacket;

  assign Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port = (1) & (Medipix_sopc_burst_7_downstream_read | Medipix_sopc_burst_7_downstream_write);
  //Medipix_sopc_burst_6/downstream granted epcs_controller/epcs_control_port last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_Medipix_sopc_burst_6_downstream_granted_slave_epcs_controller_epcs_control_port <= 0;
      else 
        last_cycle_Medipix_sopc_burst_6_downstream_granted_slave_epcs_controller_epcs_control_port <= Medipix_sopc_burst_6_downstream_saved_grant_epcs_controller_epcs_control_port ? 1 : (epcs_controller_epcs_control_port_arbitration_holdoff_internal | 0) ? 0 : last_cycle_Medipix_sopc_burst_6_downstream_granted_slave_epcs_controller_epcs_control_port;
    end


  //Medipix_sopc_burst_6_downstream_continuerequest continued request, which is an e_mux
  assign Medipix_sopc_burst_6_downstream_continuerequest = last_cycle_Medipix_sopc_burst_6_downstream_granted_slave_epcs_controller_epcs_control_port & 1;

  assign Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port = Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port & ~((Medipix_sopc_burst_7_downstream_read & ((Medipix_sopc_burst_7_downstream_latency_counter != 0))) | Medipix_sopc_burst_6_downstream_arbiterlock);
  //local readdatavalid Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port, which is an e_mux
  assign Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port = Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_7_downstream_read & ~epcs_controller_epcs_control_port_waits_for_read;

  //allow new arb cycle for epcs_controller/epcs_control_port, which is an e_assign
  assign epcs_controller_epcs_control_port_allow_new_arb_cycle = ~Medipix_sopc_burst_6_downstream_arbiterlock & ~Medipix_sopc_burst_7_downstream_arbiterlock;

  //Medipix_sopc_burst_7/downstream assignment into master qualified-requests vector for epcs_controller/epcs_control_port, which is an e_assign
  assign epcs_controller_epcs_control_port_master_qreq_vector[0] = Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port;

  //Medipix_sopc_burst_7/downstream grant epcs_controller/epcs_control_port, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port = epcs_controller_epcs_control_port_grant_vector[0];

  //Medipix_sopc_burst_7/downstream saved-grant epcs_controller/epcs_control_port, which is an e_assign
  assign Medipix_sopc_burst_7_downstream_saved_grant_epcs_controller_epcs_control_port = epcs_controller_epcs_control_port_arb_winner[0];

  //Medipix_sopc_burst_6/downstream assignment into master qualified-requests vector for epcs_controller/epcs_control_port, which is an e_assign
  assign epcs_controller_epcs_control_port_master_qreq_vector[1] = Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port;

  //Medipix_sopc_burst_6/downstream grant epcs_controller/epcs_control_port, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port = epcs_controller_epcs_control_port_grant_vector[1];

  //Medipix_sopc_burst_6/downstream saved-grant epcs_controller/epcs_control_port, which is an e_assign
  assign Medipix_sopc_burst_6_downstream_saved_grant_epcs_controller_epcs_control_port = epcs_controller_epcs_control_port_arb_winner[1];

  //epcs_controller/epcs_control_port chosen-master double-vector, which is an e_assign
  assign epcs_controller_epcs_control_port_chosen_master_double_vector = {epcs_controller_epcs_control_port_master_qreq_vector, epcs_controller_epcs_control_port_master_qreq_vector} & ({~epcs_controller_epcs_control_port_master_qreq_vector, ~epcs_controller_epcs_control_port_master_qreq_vector} + epcs_controller_epcs_control_port_arb_addend);

  //stable onehot encoding of arb winner
  assign epcs_controller_epcs_control_port_arb_winner = (epcs_controller_epcs_control_port_allow_new_arb_cycle & | epcs_controller_epcs_control_port_grant_vector) ? epcs_controller_epcs_control_port_grant_vector : epcs_controller_epcs_control_port_saved_chosen_master_vector;

  //saved epcs_controller_epcs_control_port_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_controller_epcs_control_port_saved_chosen_master_vector <= 0;
      else if (epcs_controller_epcs_control_port_allow_new_arb_cycle)
          epcs_controller_epcs_control_port_saved_chosen_master_vector <= |epcs_controller_epcs_control_port_grant_vector ? epcs_controller_epcs_control_port_grant_vector : epcs_controller_epcs_control_port_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign epcs_controller_epcs_control_port_grant_vector = {(epcs_controller_epcs_control_port_chosen_master_double_vector[1] | epcs_controller_epcs_control_port_chosen_master_double_vector[3]),
    (epcs_controller_epcs_control_port_chosen_master_double_vector[0] | epcs_controller_epcs_control_port_chosen_master_double_vector[2])};

  //epcs_controller/epcs_control_port chosen master rotated left, which is an e_assign
  assign epcs_controller_epcs_control_port_chosen_master_rot_left = (epcs_controller_epcs_control_port_arb_winner << 1) ? (epcs_controller_epcs_control_port_arb_winner << 1) : 1;

  //epcs_controller/epcs_control_port's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_controller_epcs_control_port_arb_addend <= 1;
      else if (|epcs_controller_epcs_control_port_grant_vector)
          epcs_controller_epcs_control_port_arb_addend <= epcs_controller_epcs_control_port_end_xfer? epcs_controller_epcs_control_port_chosen_master_rot_left : epcs_controller_epcs_control_port_grant_vector;
    end


  //epcs_controller_epcs_control_port_reset_n assignment, which is an e_assign
  assign epcs_controller_epcs_control_port_reset_n = reset_n;

  assign epcs_controller_epcs_control_port_chipselect = Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port | Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port;
  //epcs_controller_epcs_control_port_firsttransfer first transaction, which is an e_assign
  assign epcs_controller_epcs_control_port_firsttransfer = epcs_controller_epcs_control_port_begins_xfer ? epcs_controller_epcs_control_port_unreg_firsttransfer : epcs_controller_epcs_control_port_reg_firsttransfer;

  //epcs_controller_epcs_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign epcs_controller_epcs_control_port_unreg_firsttransfer = ~(epcs_controller_epcs_control_port_slavearbiterlockenable & epcs_controller_epcs_control_port_any_continuerequest);

  //epcs_controller_epcs_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          epcs_controller_epcs_control_port_reg_firsttransfer <= 1'b1;
      else if (epcs_controller_epcs_control_port_begins_xfer)
          epcs_controller_epcs_control_port_reg_firsttransfer <= epcs_controller_epcs_control_port_unreg_firsttransfer;
    end


  //epcs_controller_epcs_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign epcs_controller_epcs_control_port_beginbursttransfer_internal = epcs_controller_epcs_control_port_begins_xfer;

  //epcs_controller_epcs_control_port_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign epcs_controller_epcs_control_port_arbitration_holdoff_internal = epcs_controller_epcs_control_port_begins_xfer & epcs_controller_epcs_control_port_firsttransfer;

  //~epcs_controller_epcs_control_port_read_n assignment, which is an e_mux
  assign epcs_controller_epcs_control_port_read_n = ~((Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_6_downstream_read) | (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_7_downstream_read));

  //~epcs_controller_epcs_control_port_write_n assignment, which is an e_mux
  assign epcs_controller_epcs_control_port_write_n = ~((Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_6_downstream_write) | (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_7_downstream_write));

  assign shifted_address_to_epcs_controller_epcs_control_port_from_Medipix_sopc_burst_6_downstream = Medipix_sopc_burst_6_downstream_address_to_slave;
  //epcs_controller_epcs_control_port_address mux, which is an e_mux
  assign epcs_controller_epcs_control_port_address = (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port)? (shifted_address_to_epcs_controller_epcs_control_port_from_Medipix_sopc_burst_6_downstream >> 2) :
    (shifted_address_to_epcs_controller_epcs_control_port_from_Medipix_sopc_burst_7_downstream >> 2);

  assign shifted_address_to_epcs_controller_epcs_control_port_from_Medipix_sopc_burst_7_downstream = Medipix_sopc_burst_7_downstream_address_to_slave;
  //d1_epcs_controller_epcs_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_epcs_controller_epcs_control_port_end_xfer <= 1;
      else 
        d1_epcs_controller_epcs_control_port_end_xfer <= epcs_controller_epcs_control_port_end_xfer;
    end


  //epcs_controller_epcs_control_port_waits_for_read in a cycle, which is an e_mux
  assign epcs_controller_epcs_control_port_waits_for_read = epcs_controller_epcs_control_port_in_a_read_cycle & epcs_controller_epcs_control_port_begins_xfer;

  //epcs_controller_epcs_control_port_in_a_read_cycle assignment, which is an e_assign
  assign epcs_controller_epcs_control_port_in_a_read_cycle = (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_6_downstream_read) | (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_7_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = epcs_controller_epcs_control_port_in_a_read_cycle;

  //epcs_controller_epcs_control_port_waits_for_write in a cycle, which is an e_mux
  assign epcs_controller_epcs_control_port_waits_for_write = epcs_controller_epcs_control_port_in_a_write_cycle & epcs_controller_epcs_control_port_begins_xfer;

  //epcs_controller_epcs_control_port_in_a_write_cycle assignment, which is an e_assign
  assign epcs_controller_epcs_control_port_in_a_write_cycle = (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_6_downstream_write) | (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port & Medipix_sopc_burst_7_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = epcs_controller_epcs_control_port_in_a_write_cycle;

  assign wait_for_epcs_controller_epcs_control_port_counter = 0;
  //assign epcs_controller_epcs_control_port_irq_from_sa = epcs_controller_epcs_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign epcs_controller_epcs_control_port_irq_from_sa = epcs_controller_epcs_control_port_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //epcs_controller/epcs_control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_6/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port && (Medipix_sopc_burst_6_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_6/downstream drove 0 on its 'arbitrationshare' port while accessing slave epcs_controller/epcs_control_port", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_6/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port && (Medipix_sopc_burst_6_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_6/downstream drove 0 on its 'burstcount' port while accessing slave epcs_controller/epcs_control_port", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port && (Medipix_sopc_burst_7_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_7/downstream drove 0 on its 'arbitrationshare' port while accessing slave epcs_controller/epcs_control_port", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_7/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port && (Medipix_sopc_burst_7_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_7/downstream drove 0 on its 'burstcount' port while accessing slave epcs_controller/epcs_control_port", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port + Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_6_downstream_saved_grant_epcs_controller_epcs_control_port + Medipix_sopc_burst_7_downstream_saved_grant_epcs_controller_epcs_control_port > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module igor_mac_control_port_arbitrator (
                                          // inputs:
                                           Medipix_sopc_burst_8_downstream_address_to_slave,
                                           Medipix_sopc_burst_8_downstream_arbitrationshare,
                                           Medipix_sopc_burst_8_downstream_burstcount,
                                           Medipix_sopc_burst_8_downstream_latency_counter,
                                           Medipix_sopc_burst_8_downstream_read,
                                           Medipix_sopc_burst_8_downstream_write,
                                           Medipix_sopc_burst_8_downstream_writedata,
                                           clk,
                                           igor_mac_control_port_irq,
                                           igor_mac_control_port_readdata,
                                           igor_mac_control_port_waitrequest_n,
                                           reset_n,

                                          // outputs:
                                           Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port,
                                           Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port,
                                           Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port,
                                           Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port,
                                           d1_igor_mac_control_port_end_xfer,
                                           igor_mac_control_port_address,
                                           igor_mac_control_port_chipselect,
                                           igor_mac_control_port_irq_from_sa,
                                           igor_mac_control_port_read,
                                           igor_mac_control_port_readdata_from_sa,
                                           igor_mac_control_port_reset,
                                           igor_mac_control_port_waitrequest_n_from_sa,
                                           igor_mac_control_port_write,
                                           igor_mac_control_port_writedata
                                        )
;

  output           Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port;
  output           Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port;
  output           Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port;
  output           Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port;
  output           d1_igor_mac_control_port_end_xfer;
  output  [  9: 0] igor_mac_control_port_address;
  output           igor_mac_control_port_chipselect;
  output           igor_mac_control_port_irq_from_sa;
  output           igor_mac_control_port_read;
  output  [ 31: 0] igor_mac_control_port_readdata_from_sa;
  output           igor_mac_control_port_reset;
  output           igor_mac_control_port_waitrequest_n_from_sa;
  output           igor_mac_control_port_write;
  output  [ 31: 0] igor_mac_control_port_writedata;
  input   [ 11: 0] Medipix_sopc_burst_8_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_8_downstream_arbitrationshare;
  input            Medipix_sopc_burst_8_downstream_burstcount;
  input            Medipix_sopc_burst_8_downstream_latency_counter;
  input            Medipix_sopc_burst_8_downstream_read;
  input            Medipix_sopc_burst_8_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_8_downstream_writedata;
  input            clk;
  input            igor_mac_control_port_irq;
  input   [ 31: 0] igor_mac_control_port_readdata;
  input            igor_mac_control_port_waitrequest_n;
  input            reset_n;

  wire             Medipix_sopc_burst_8_downstream_arbiterlock;
  wire             Medipix_sopc_burst_8_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_8_downstream_continuerequest;
  wire             Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_saved_grant_igor_mac_control_port;
  reg              d1_igor_mac_control_port_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_igor_mac_control_port;
  wire    [  9: 0] igor_mac_control_port_address;
  wire             igor_mac_control_port_allgrants;
  wire             igor_mac_control_port_allow_new_arb_cycle;
  wire             igor_mac_control_port_any_bursting_master_saved_grant;
  wire             igor_mac_control_port_any_continuerequest;
  wire             igor_mac_control_port_arb_counter_enable;
  reg     [  3: 0] igor_mac_control_port_arb_share_counter;
  wire    [  3: 0] igor_mac_control_port_arb_share_counter_next_value;
  wire    [  3: 0] igor_mac_control_port_arb_share_set_values;
  wire             igor_mac_control_port_beginbursttransfer_internal;
  wire             igor_mac_control_port_begins_xfer;
  wire             igor_mac_control_port_chipselect;
  wire             igor_mac_control_port_end_xfer;
  wire             igor_mac_control_port_firsttransfer;
  wire             igor_mac_control_port_grant_vector;
  wire             igor_mac_control_port_in_a_read_cycle;
  wire             igor_mac_control_port_in_a_write_cycle;
  wire             igor_mac_control_port_irq_from_sa;
  wire             igor_mac_control_port_master_qreq_vector;
  wire             igor_mac_control_port_non_bursting_master_requests;
  wire             igor_mac_control_port_read;
  wire    [ 31: 0] igor_mac_control_port_readdata_from_sa;
  reg              igor_mac_control_port_reg_firsttransfer;
  wire             igor_mac_control_port_reset;
  reg              igor_mac_control_port_slavearbiterlockenable;
  wire             igor_mac_control_port_slavearbiterlockenable2;
  wire             igor_mac_control_port_unreg_firsttransfer;
  wire             igor_mac_control_port_waitrequest_n_from_sa;
  wire             igor_mac_control_port_waits_for_read;
  wire             igor_mac_control_port_waits_for_write;
  wire             igor_mac_control_port_write;
  wire    [ 31: 0] igor_mac_control_port_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 11: 0] shifted_address_to_igor_mac_control_port_from_Medipix_sopc_burst_8_downstream;
  wire             wait_for_igor_mac_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~igor_mac_control_port_end_xfer;
    end


  assign igor_mac_control_port_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port));
  //assign igor_mac_control_port_readdata_from_sa = igor_mac_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign igor_mac_control_port_readdata_from_sa = igor_mac_control_port_readdata;

  assign Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port = (1) & (Medipix_sopc_burst_8_downstream_read | Medipix_sopc_burst_8_downstream_write);
  //assign igor_mac_control_port_waitrequest_n_from_sa = igor_mac_control_port_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign igor_mac_control_port_waitrequest_n_from_sa = igor_mac_control_port_waitrequest_n;

  //igor_mac_control_port_arb_share_counter set values, which is an e_mux
  assign igor_mac_control_port_arb_share_set_values = (Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port)? Medipix_sopc_burst_8_downstream_arbitrationshare :
    1;

  //igor_mac_control_port_non_bursting_master_requests mux, which is an e_mux
  assign igor_mac_control_port_non_bursting_master_requests = 0;

  //igor_mac_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign igor_mac_control_port_any_bursting_master_saved_grant = Medipix_sopc_burst_8_downstream_saved_grant_igor_mac_control_port;

  //igor_mac_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign igor_mac_control_port_arb_share_counter_next_value = igor_mac_control_port_firsttransfer ? (igor_mac_control_port_arb_share_set_values - 1) : |igor_mac_control_port_arb_share_counter ? (igor_mac_control_port_arb_share_counter - 1) : 0;

  //igor_mac_control_port_allgrants all slave grants, which is an e_mux
  assign igor_mac_control_port_allgrants = |igor_mac_control_port_grant_vector;

  //igor_mac_control_port_end_xfer assignment, which is an e_assign
  assign igor_mac_control_port_end_xfer = ~(igor_mac_control_port_waits_for_read | igor_mac_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_igor_mac_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_igor_mac_control_port = igor_mac_control_port_end_xfer & (~igor_mac_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //igor_mac_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign igor_mac_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_igor_mac_control_port & igor_mac_control_port_allgrants) | (end_xfer_arb_share_counter_term_igor_mac_control_port & ~igor_mac_control_port_non_bursting_master_requests);

  //igor_mac_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_control_port_arb_share_counter <= 0;
      else if (igor_mac_control_port_arb_counter_enable)
          igor_mac_control_port_arb_share_counter <= igor_mac_control_port_arb_share_counter_next_value;
    end


  //igor_mac_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_control_port_slavearbiterlockenable <= 0;
      else if ((|igor_mac_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_igor_mac_control_port) | (end_xfer_arb_share_counter_term_igor_mac_control_port & ~igor_mac_control_port_non_bursting_master_requests))
          igor_mac_control_port_slavearbiterlockenable <= |igor_mac_control_port_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_8/downstream igor_mac/control_port arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_arbiterlock = igor_mac_control_port_slavearbiterlockenable & Medipix_sopc_burst_8_downstream_continuerequest;

  //igor_mac_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign igor_mac_control_port_slavearbiterlockenable2 = |igor_mac_control_port_arb_share_counter_next_value;

  //Medipix_sopc_burst_8/downstream igor_mac/control_port arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_arbiterlock2 = igor_mac_control_port_slavearbiterlockenable2 & Medipix_sopc_burst_8_downstream_continuerequest;

  //igor_mac_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  assign igor_mac_control_port_any_continuerequest = 1;

  //Medipix_sopc_burst_8_downstream_continuerequest continued request, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_continuerequest = 1;

  assign Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port = Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port & ~((Medipix_sopc_burst_8_downstream_read & ((Medipix_sopc_burst_8_downstream_latency_counter != 0))));
  //local readdatavalid Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port, which is an e_mux
  assign Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port = Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port & Medipix_sopc_burst_8_downstream_read & ~igor_mac_control_port_waits_for_read;

  //igor_mac_control_port_writedata mux, which is an e_mux
  assign igor_mac_control_port_writedata = Medipix_sopc_burst_8_downstream_writedata;

  //master is always granted when requested
  assign Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port = Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port;

  //Medipix_sopc_burst_8/downstream saved-grant igor_mac/control_port, which is an e_assign
  assign Medipix_sopc_burst_8_downstream_saved_grant_igor_mac_control_port = Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port;

  //allow new arb cycle for igor_mac/control_port, which is an e_assign
  assign igor_mac_control_port_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign igor_mac_control_port_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign igor_mac_control_port_master_qreq_vector = 1;

  //~igor_mac_control_port_reset assignment, which is an e_assign
  assign igor_mac_control_port_reset = ~reset_n;

  assign igor_mac_control_port_chipselect = Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port;
  //igor_mac_control_port_firsttransfer first transaction, which is an e_assign
  assign igor_mac_control_port_firsttransfer = igor_mac_control_port_begins_xfer ? igor_mac_control_port_unreg_firsttransfer : igor_mac_control_port_reg_firsttransfer;

  //igor_mac_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign igor_mac_control_port_unreg_firsttransfer = ~(igor_mac_control_port_slavearbiterlockenable & igor_mac_control_port_any_continuerequest);

  //igor_mac_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_control_port_reg_firsttransfer <= 1'b1;
      else if (igor_mac_control_port_begins_xfer)
          igor_mac_control_port_reg_firsttransfer <= igor_mac_control_port_unreg_firsttransfer;
    end


  //igor_mac_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign igor_mac_control_port_beginbursttransfer_internal = igor_mac_control_port_begins_xfer;

  //igor_mac_control_port_read assignment, which is an e_mux
  assign igor_mac_control_port_read = Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port & Medipix_sopc_burst_8_downstream_read;

  //igor_mac_control_port_write assignment, which is an e_mux
  assign igor_mac_control_port_write = Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port & Medipix_sopc_burst_8_downstream_write;

  assign shifted_address_to_igor_mac_control_port_from_Medipix_sopc_burst_8_downstream = Medipix_sopc_burst_8_downstream_address_to_slave;
  //igor_mac_control_port_address mux, which is an e_mux
  assign igor_mac_control_port_address = shifted_address_to_igor_mac_control_port_from_Medipix_sopc_burst_8_downstream >> 2;

  //d1_igor_mac_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_igor_mac_control_port_end_xfer <= 1;
      else 
        d1_igor_mac_control_port_end_xfer <= igor_mac_control_port_end_xfer;
    end


  //igor_mac_control_port_waits_for_read in a cycle, which is an e_mux
  assign igor_mac_control_port_waits_for_read = igor_mac_control_port_in_a_read_cycle & ~igor_mac_control_port_waitrequest_n_from_sa;

  //igor_mac_control_port_in_a_read_cycle assignment, which is an e_assign
  assign igor_mac_control_port_in_a_read_cycle = Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port & Medipix_sopc_burst_8_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = igor_mac_control_port_in_a_read_cycle;

  //igor_mac_control_port_waits_for_write in a cycle, which is an e_mux
  assign igor_mac_control_port_waits_for_write = igor_mac_control_port_in_a_write_cycle & ~igor_mac_control_port_waitrequest_n_from_sa;

  //igor_mac_control_port_in_a_write_cycle assignment, which is an e_assign
  assign igor_mac_control_port_in_a_write_cycle = Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port & Medipix_sopc_burst_8_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = igor_mac_control_port_in_a_write_cycle;

  assign wait_for_igor_mac_control_port_counter = 0;
  //assign igor_mac_control_port_irq_from_sa = igor_mac_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign igor_mac_control_port_irq_from_sa = igor_mac_control_port_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //igor_mac/control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_8/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port && (Medipix_sopc_burst_8_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_8/downstream drove 0 on its 'arbitrationshare' port while accessing slave igor_mac/control_port", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_8/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port && (Medipix_sopc_burst_8_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_8/downstream drove 0 on its 'burstcount' port while accessing slave igor_mac/control_port", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module igor_mac_rx_master_arbitrator (
                                       // inputs:
                                        clk,
                                        clock_crossing_s1_waitrequest_from_sa,
                                        d1_clock_crossing_s1_end_xfer,
                                        igor_mac_rx_master_address,
                                        igor_mac_rx_master_byteenable,
                                        igor_mac_rx_master_granted_clock_crossing_s1,
                                        igor_mac_rx_master_qualified_request_clock_crossing_s1,
                                        igor_mac_rx_master_requests_clock_crossing_s1,
                                        igor_mac_rx_master_write,
                                        igor_mac_rx_master_writedata,
                                        reset_n,

                                       // outputs:
                                        igor_mac_rx_master_address_to_slave,
                                        igor_mac_rx_master_waitrequest
                                     )
;

  output  [ 31: 0] igor_mac_rx_master_address_to_slave;
  output           igor_mac_rx_master_waitrequest;
  input            clk;
  input            clock_crossing_s1_waitrequest_from_sa;
  input            d1_clock_crossing_s1_end_xfer;
  input   [ 31: 0] igor_mac_rx_master_address;
  input   [  3: 0] igor_mac_rx_master_byteenable;
  input            igor_mac_rx_master_granted_clock_crossing_s1;
  input            igor_mac_rx_master_qualified_request_clock_crossing_s1;
  input            igor_mac_rx_master_requests_clock_crossing_s1;
  input            igor_mac_rx_master_write;
  input   [ 31: 0] igor_mac_rx_master_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 31: 0] igor_mac_rx_master_address_last_time;
  wire    [ 31: 0] igor_mac_rx_master_address_to_slave;
  reg     [  3: 0] igor_mac_rx_master_byteenable_last_time;
  wire             igor_mac_rx_master_run;
  wire             igor_mac_rx_master_waitrequest;
  reg              igor_mac_rx_master_write_last_time;
  reg     [ 31: 0] igor_mac_rx_master_writedata_last_time;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (igor_mac_rx_master_qualified_request_clock_crossing_s1 | ~igor_mac_rx_master_requests_clock_crossing_s1) & (igor_mac_rx_master_granted_clock_crossing_s1 | ~igor_mac_rx_master_qualified_request_clock_crossing_s1) & ((~igor_mac_rx_master_qualified_request_clock_crossing_s1 | ~(igor_mac_rx_master_write) | (1 & ~clock_crossing_s1_waitrequest_from_sa & (igor_mac_rx_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign igor_mac_rx_master_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign igor_mac_rx_master_address_to_slave = {5'b0,
    igor_mac_rx_master_address[26 : 0]};

  //actual waitrequest port, which is an e_assign
  assign igor_mac_rx_master_waitrequest = ~igor_mac_rx_master_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //igor_mac_rx_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_rx_master_address_last_time <= 0;
      else 
        igor_mac_rx_master_address_last_time <= igor_mac_rx_master_address;
    end


  //igor_mac/rx_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= igor_mac_rx_master_waitrequest & (igor_mac_rx_master_write);
    end


  //igor_mac_rx_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (igor_mac_rx_master_address != igor_mac_rx_master_address_last_time))
        begin
          $write("%0d ns: igor_mac_rx_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //igor_mac_rx_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_rx_master_byteenable_last_time <= 0;
      else 
        igor_mac_rx_master_byteenable_last_time <= igor_mac_rx_master_byteenable;
    end


  //igor_mac_rx_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (igor_mac_rx_master_byteenable != igor_mac_rx_master_byteenable_last_time))
        begin
          $write("%0d ns: igor_mac_rx_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //igor_mac_rx_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_rx_master_write_last_time <= 0;
      else 
        igor_mac_rx_master_write_last_time <= igor_mac_rx_master_write;
    end


  //igor_mac_rx_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (igor_mac_rx_master_write != igor_mac_rx_master_write_last_time))
        begin
          $write("%0d ns: igor_mac_rx_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //igor_mac_rx_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_rx_master_writedata_last_time <= 0;
      else 
        igor_mac_rx_master_writedata_last_time <= igor_mac_rx_master_writedata;
    end


  //igor_mac_rx_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (igor_mac_rx_master_writedata != igor_mac_rx_master_writedata_last_time) & igor_mac_rx_master_write)
        begin
          $write("%0d ns: igor_mac_rx_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module igor_mac_tx_master_arbitrator (
                                       // inputs:
                                        clk,
                                        clock_crossing_s1_readdata_from_sa,
                                        clock_crossing_s1_waitrequest_from_sa,
                                        d1_clock_crossing_s1_end_xfer,
                                        igor_mac_tx_master_address,
                                        igor_mac_tx_master_granted_clock_crossing_s1,
                                        igor_mac_tx_master_qualified_request_clock_crossing_s1,
                                        igor_mac_tx_master_read,
                                        igor_mac_tx_master_read_data_valid_clock_crossing_s1,
                                        igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register,
                                        igor_mac_tx_master_requests_clock_crossing_s1,
                                        reset_n,

                                       // outputs:
                                        igor_mac_tx_master_address_to_slave,
                                        igor_mac_tx_master_latency_counter,
                                        igor_mac_tx_master_readdata,
                                        igor_mac_tx_master_readdatavalid,
                                        igor_mac_tx_master_waitrequest
                                     )
;

  output  [ 31: 0] igor_mac_tx_master_address_to_slave;
  output           igor_mac_tx_master_latency_counter;
  output  [ 31: 0] igor_mac_tx_master_readdata;
  output           igor_mac_tx_master_readdatavalid;
  output           igor_mac_tx_master_waitrequest;
  input            clk;
  input   [ 31: 0] clock_crossing_s1_readdata_from_sa;
  input            clock_crossing_s1_waitrequest_from_sa;
  input            d1_clock_crossing_s1_end_xfer;
  input   [ 31: 0] igor_mac_tx_master_address;
  input            igor_mac_tx_master_granted_clock_crossing_s1;
  input            igor_mac_tx_master_qualified_request_clock_crossing_s1;
  input            igor_mac_tx_master_read;
  input            igor_mac_tx_master_read_data_valid_clock_crossing_s1;
  input            igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register;
  input            igor_mac_tx_master_requests_clock_crossing_s1;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 31: 0] igor_mac_tx_master_address_last_time;
  wire    [ 31: 0] igor_mac_tx_master_address_to_slave;
  wire             igor_mac_tx_master_is_granted_some_slave;
  reg              igor_mac_tx_master_latency_counter;
  reg              igor_mac_tx_master_read_but_no_slave_selected;
  reg              igor_mac_tx_master_read_last_time;
  wire    [ 31: 0] igor_mac_tx_master_readdata;
  wire             igor_mac_tx_master_readdatavalid;
  wire             igor_mac_tx_master_run;
  wire             igor_mac_tx_master_waitrequest;
  wire             latency_load_value;
  wire             p1_igor_mac_tx_master_latency_counter;
  wire             pre_flush_igor_mac_tx_master_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (igor_mac_tx_master_qualified_request_clock_crossing_s1 | ~igor_mac_tx_master_requests_clock_crossing_s1) & (igor_mac_tx_master_granted_clock_crossing_s1 | ~igor_mac_tx_master_qualified_request_clock_crossing_s1) & ((~igor_mac_tx_master_qualified_request_clock_crossing_s1 | ~(igor_mac_tx_master_read) | (1 & ~clock_crossing_s1_waitrequest_from_sa & (igor_mac_tx_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign igor_mac_tx_master_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign igor_mac_tx_master_address_to_slave = {5'b0,
    igor_mac_tx_master_address[26 : 0]};

  //igor_mac_tx_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_tx_master_read_but_no_slave_selected <= 0;
      else 
        igor_mac_tx_master_read_but_no_slave_selected <= igor_mac_tx_master_read & igor_mac_tx_master_run & ~igor_mac_tx_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign igor_mac_tx_master_is_granted_some_slave = igor_mac_tx_master_granted_clock_crossing_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_igor_mac_tx_master_readdatavalid = igor_mac_tx_master_read_data_valid_clock_crossing_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign igor_mac_tx_master_readdatavalid = igor_mac_tx_master_read_but_no_slave_selected |
    pre_flush_igor_mac_tx_master_readdatavalid;

  //igor_mac/tx_master readdata mux, which is an e_mux
  assign igor_mac_tx_master_readdata = clock_crossing_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign igor_mac_tx_master_waitrequest = ~igor_mac_tx_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_tx_master_latency_counter <= 0;
      else 
        igor_mac_tx_master_latency_counter <= p1_igor_mac_tx_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_igor_mac_tx_master_latency_counter = ((igor_mac_tx_master_run & igor_mac_tx_master_read))? latency_load_value :
    (igor_mac_tx_master_latency_counter)? igor_mac_tx_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //igor_mac_tx_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_tx_master_address_last_time <= 0;
      else 
        igor_mac_tx_master_address_last_time <= igor_mac_tx_master_address;
    end


  //igor_mac/tx_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= igor_mac_tx_master_waitrequest & (igor_mac_tx_master_read);
    end


  //igor_mac_tx_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (igor_mac_tx_master_address != igor_mac_tx_master_address_last_time))
        begin
          $write("%0d ns: igor_mac_tx_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //igor_mac_tx_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          igor_mac_tx_master_read_last_time <= 0;
      else 
        igor_mac_tx_master_read_last_time <= igor_mac_tx_master_read;
    end


  //igor_mac_tx_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (igor_mac_tx_master_read != igor_mac_tx_master_read_last_time))
        begin
          $write("%0d ns: igor_mac_tx_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_0_avalon_jtag_slave_arbitrator (
                                                  // inputs:
                                                   Medipix_sopc_burst_2_downstream_address_to_slave,
                                                   Medipix_sopc_burst_2_downstream_arbitrationshare,
                                                   Medipix_sopc_burst_2_downstream_burstcount,
                                                   Medipix_sopc_burst_2_downstream_latency_counter,
                                                   Medipix_sopc_burst_2_downstream_nativeaddress,
                                                   Medipix_sopc_burst_2_downstream_read,
                                                   Medipix_sopc_burst_2_downstream_write,
                                                   Medipix_sopc_burst_2_downstream_writedata,
                                                   clk,
                                                   jtag_uart_0_avalon_jtag_slave_dataavailable,
                                                   jtag_uart_0_avalon_jtag_slave_irq,
                                                   jtag_uart_0_avalon_jtag_slave_readdata,
                                                   jtag_uart_0_avalon_jtag_slave_readyfordata,
                                                   jtag_uart_0_avalon_jtag_slave_waitrequest,
                                                   reset_n,

                                                  // outputs:
                                                   Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave,
                                                   Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave,
                                                   Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave,
                                                   Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave,
                                                   d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
                                                   jtag_uart_0_avalon_jtag_slave_address,
                                                   jtag_uart_0_avalon_jtag_slave_chipselect,
                                                   jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_irq_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_read_n,
                                                   jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_reset_n,
                                                   jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_write_n,
                                                   jtag_uart_0_avalon_jtag_slave_writedata
                                                )
;

  output           Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave;
  output           Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave;
  output           Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  output           Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave;
  output           d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  output           jtag_uart_0_avalon_jtag_slave_address;
  output           jtag_uart_0_avalon_jtag_slave_chipselect;
  output           jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_reset_n;
  output           jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  input   [  2: 0] Medipix_sopc_burst_2_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_2_downstream_arbitrationshare;
  input            Medipix_sopc_burst_2_downstream_burstcount;
  input            Medipix_sopc_burst_2_downstream_latency_counter;
  input   [  2: 0] Medipix_sopc_burst_2_downstream_nativeaddress;
  input            Medipix_sopc_burst_2_downstream_read;
  input            Medipix_sopc_burst_2_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_2_downstream_writedata;
  input            clk;
  input            jtag_uart_0_avalon_jtag_slave_dataavailable;
  input            jtag_uart_0_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata;
  input            jtag_uart_0_avalon_jtag_slave_readyfordata;
  input            jtag_uart_0_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             Medipix_sopc_burst_2_downstream_arbiterlock;
  wire             Medipix_sopc_burst_2_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_2_downstream_continuerequest;
  wire             Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_saved_grant_jtag_uart_0_avalon_jtag_slave;
  reg              d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_address;
  wire             jtag_uart_0_avalon_jtag_slave_allgrants;
  wire             jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_0_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_0_avalon_jtag_slave_arb_counter_enable;
  reg     [  3: 0] jtag_uart_0_avalon_jtag_slave_arb_share_counter;
  wire    [  3: 0] jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  3: 0] jtag_uart_0_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_0_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_chipselect;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_0_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_0_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_reset_n;
  reg              jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_0_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_0_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  wire             wait_for_jtag_uart_0_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_0_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_0_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave));
  //assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata;

  assign Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave = (1) & (Medipix_sopc_burst_2_downstream_read | Medipix_sopc_burst_2_downstream_write);
  //assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest;

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_arb_share_set_values = (Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave)? Medipix_sopc_burst_2_downstream_arbitrationshare :
    1;

  //jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests = 0;

  //jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant = Medipix_sopc_burst_2_downstream_saved_grant_jtag_uart_0_avalon_jtag_slave;

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_0_avalon_jtag_slave_firsttransfer ? (jtag_uart_0_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_0_avalon_jtag_slave_arb_share_counter ? (jtag_uart_0_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_0_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_allgrants = |jtag_uart_0_avalon_jtag_slave_grant_vector;

  //jtag_uart_0_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_end_xfer = ~(jtag_uart_0_avalon_jtag_slave_waits_for_read | jtag_uart_0_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave = jtag_uart_0_avalon_jtag_slave_end_xfer & (~jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & jtag_uart_0_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & ~jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_0_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_0_avalon_jtag_slave_arb_share_counter <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_0_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & ~jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_2/downstream jtag_uart_0/avalon_jtag_slave arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_arbiterlock = jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable & Medipix_sopc_burst_2_downstream_continuerequest;

  //jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;

  //Medipix_sopc_burst_2/downstream jtag_uart_0/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_arbiterlock2 = jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 & Medipix_sopc_burst_2_downstream_continuerequest;

  //jtag_uart_0_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_any_continuerequest = 1;

  //Medipix_sopc_burst_2_downstream_continuerequest continued request, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_continuerequest = 1;

  assign Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave = Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave & ~((Medipix_sopc_burst_2_downstream_read & ((Medipix_sopc_burst_2_downstream_latency_counter != 0))));
  //local readdatavalid Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave, which is an e_mux
  assign Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave = Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave & Medipix_sopc_burst_2_downstream_read & ~jtag_uart_0_avalon_jtag_slave_waits_for_read;

  //jtag_uart_0_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_writedata = Medipix_sopc_burst_2_downstream_writedata;

  //master is always granted when requested
  assign Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave = Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave;

  //Medipix_sopc_burst_2/downstream saved-grant jtag_uart_0/avalon_jtag_slave, which is an e_assign
  assign Medipix_sopc_burst_2_downstream_saved_grant_jtag_uart_0_avalon_jtag_slave = Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart_0/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_0_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_0_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_0_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_0_avalon_jtag_slave_chipselect = Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave;
  //jtag_uart_0_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_firsttransfer = jtag_uart_0_avalon_jtag_slave_begins_xfer ? jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_0_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_0_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_0_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_0_avalon_jtag_slave_begins_xfer)
          jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_0_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_0_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_read_n = ~(Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave & Medipix_sopc_burst_2_downstream_read);

  //~jtag_uart_0_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_write_n = ~(Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave & Medipix_sopc_burst_2_downstream_write);

  //jtag_uart_0_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_address = Medipix_sopc_burst_2_downstream_nativeaddress;

  //d1_jtag_uart_0_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= jtag_uart_0_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_0_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_waits_for_read = jtag_uart_0_avalon_jtag_slave_in_a_read_cycle & jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_0_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_in_a_read_cycle = Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave & Medipix_sopc_burst_2_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_0_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_waits_for_write = jtag_uart_0_avalon_jtag_slave_in_a_write_cycle & jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_0_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_in_a_write_cycle = Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave & Medipix_sopc_burst_2_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_0_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_0/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_2/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave && (Medipix_sopc_burst_2_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_2/downstream drove 0 on its 'arbitrationshare' port while accessing slave jtag_uart_0/avalon_jtag_slave", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_2/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave && (Medipix_sopc_burst_2_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_2/downstream drove 0 on its 'burstcount' port while accessing slave jtag_uart_0/avalon_jtag_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_clock_crossing_m1_to_ram_s1_module (
                                                         // inputs:
                                                          clear_fifo,
                                                          clk,
                                                          data_in,
                                                          read,
                                                          reset_n,
                                                          sync_reset,
                                                          write,

                                                         // outputs:
                                                          data_out,
                                                          empty,
                                                          fifo_contains_ones_n,
                                                          full
                                                       )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ram_s1_arbitrator (
                           // inputs:
                            clk,
                            clock_crossing_m1_address_to_slave,
                            clock_crossing_m1_byteenable,
                            clock_crossing_m1_latency_counter,
                            clock_crossing_m1_read,
                            clock_crossing_m1_write,
                            clock_crossing_m1_writedata,
                            ram_s1_readdata,
                            ram_s1_readdatavalid,
                            ram_s1_resetrequest_n,
                            ram_s1_waitrequest_n,
                            reset_n,

                           // outputs:
                            clock_crossing_m1_granted_ram_s1,
                            clock_crossing_m1_qualified_request_ram_s1,
                            clock_crossing_m1_read_data_valid_ram_s1,
                            clock_crossing_m1_read_data_valid_ram_s1_shift_register,
                            clock_crossing_m1_requests_ram_s1,
                            d1_ram_s1_end_xfer,
                            ram_s1_address,
                            ram_s1_beginbursttransfer,
                            ram_s1_burstcount,
                            ram_s1_byteenable,
                            ram_s1_read,
                            ram_s1_readdata_from_sa,
                            ram_s1_resetrequest_n_from_sa,
                            ram_s1_waitrequest_n_from_sa,
                            ram_s1_write,
                            ram_s1_writedata
                         )
;

  output           clock_crossing_m1_granted_ram_s1;
  output           clock_crossing_m1_qualified_request_ram_s1;
  output           clock_crossing_m1_read_data_valid_ram_s1;
  output           clock_crossing_m1_read_data_valid_ram_s1_shift_register;
  output           clock_crossing_m1_requests_ram_s1;
  output           d1_ram_s1_end_xfer;
  output  [ 24: 0] ram_s1_address;
  output           ram_s1_beginbursttransfer;
  output  [  2: 0] ram_s1_burstcount;
  output  [  3: 0] ram_s1_byteenable;
  output           ram_s1_read;
  output  [ 31: 0] ram_s1_readdata_from_sa;
  output           ram_s1_resetrequest_n_from_sa;
  output           ram_s1_waitrequest_n_from_sa;
  output           ram_s1_write;
  output  [ 31: 0] ram_s1_writedata;
  input            clk;
  input   [ 26: 0] clock_crossing_m1_address_to_slave;
  input   [  3: 0] clock_crossing_m1_byteenable;
  input            clock_crossing_m1_latency_counter;
  input            clock_crossing_m1_read;
  input            clock_crossing_m1_write;
  input   [ 31: 0] clock_crossing_m1_writedata;
  input   [ 31: 0] ram_s1_readdata;
  input            ram_s1_readdatavalid;
  input            ram_s1_resetrequest_n;
  input            ram_s1_waitrequest_n;
  input            reset_n;

  wire             clock_crossing_m1_arbiterlock;
  wire             clock_crossing_m1_arbiterlock2;
  wire             clock_crossing_m1_continuerequest;
  wire             clock_crossing_m1_granted_ram_s1;
  wire             clock_crossing_m1_qualified_request_ram_s1;
  wire             clock_crossing_m1_rdv_fifo_empty_ram_s1;
  wire             clock_crossing_m1_rdv_fifo_output_from_ram_s1;
  wire             clock_crossing_m1_read_data_valid_ram_s1;
  wire             clock_crossing_m1_read_data_valid_ram_s1_shift_register;
  wire             clock_crossing_m1_requests_ram_s1;
  wire             clock_crossing_m1_saved_grant_ram_s1;
  reg              d1_ram_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 24: 0] ram_s1_address;
  wire             ram_s1_allgrants;
  wire             ram_s1_allow_new_arb_cycle;
  wire             ram_s1_any_bursting_master_saved_grant;
  wire             ram_s1_any_continuerequest;
  wire             ram_s1_arb_counter_enable;
  reg              ram_s1_arb_share_counter;
  wire             ram_s1_arb_share_counter_next_value;
  wire             ram_s1_arb_share_set_values;
  reg     [  1: 0] ram_s1_bbt_burstcounter;
  wire             ram_s1_beginbursttransfer;
  wire             ram_s1_beginbursttransfer_internal;
  wire             ram_s1_begins_xfer;
  wire    [  2: 0] ram_s1_burstcount;
  wire    [  3: 0] ram_s1_byteenable;
  wire             ram_s1_end_xfer;
  wire             ram_s1_firsttransfer;
  wire             ram_s1_grant_vector;
  wire             ram_s1_in_a_read_cycle;
  wire             ram_s1_in_a_write_cycle;
  wire             ram_s1_master_qreq_vector;
  wire             ram_s1_move_on_to_next_transaction;
  wire    [  1: 0] ram_s1_next_bbt_burstcount;
  wire             ram_s1_non_bursting_master_requests;
  wire             ram_s1_read;
  wire    [ 31: 0] ram_s1_readdata_from_sa;
  wire             ram_s1_readdatavalid_from_sa;
  reg              ram_s1_reg_firsttransfer;
  wire             ram_s1_resetrequest_n_from_sa;
  reg              ram_s1_slavearbiterlockenable;
  wire             ram_s1_slavearbiterlockenable2;
  wire             ram_s1_unreg_firsttransfer;
  wire             ram_s1_waitrequest_n_from_sa;
  wire             ram_s1_waits_for_read;
  wire             ram_s1_waits_for_write;
  wire             ram_s1_write;
  wire    [ 31: 0] ram_s1_writedata;
  wire    [ 26: 0] shifted_address_to_ram_s1_from_clock_crossing_m1;
  wire             wait_for_ram_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ram_s1_end_xfer;
    end


  assign ram_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_m1_qualified_request_ram_s1));
  //assign ram_s1_readdata_from_sa = ram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ram_s1_readdata_from_sa = ram_s1_readdata;

  assign clock_crossing_m1_requests_ram_s1 = (1) & (clock_crossing_m1_read | clock_crossing_m1_write);
  //assign ram_s1_waitrequest_n_from_sa = ram_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ram_s1_waitrequest_n_from_sa = ram_s1_waitrequest_n;

  //assign ram_s1_readdatavalid_from_sa = ram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ram_s1_readdatavalid_from_sa = ram_s1_readdatavalid;

  //ram_s1_arb_share_counter set values, which is an e_mux
  assign ram_s1_arb_share_set_values = 1;

  //ram_s1_non_bursting_master_requests mux, which is an e_mux
  assign ram_s1_non_bursting_master_requests = clock_crossing_m1_requests_ram_s1;

  //ram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ram_s1_any_bursting_master_saved_grant = 0;

  //ram_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ram_s1_arb_share_counter_next_value = ram_s1_firsttransfer ? (ram_s1_arb_share_set_values - 1) : |ram_s1_arb_share_counter ? (ram_s1_arb_share_counter - 1) : 0;

  //ram_s1_allgrants all slave grants, which is an e_mux
  assign ram_s1_allgrants = |ram_s1_grant_vector;

  //ram_s1_end_xfer assignment, which is an e_assign
  assign ram_s1_end_xfer = ~(ram_s1_waits_for_read | ram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ram_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ram_s1 = ram_s1_end_xfer & (~ram_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ram_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ram_s1 & ram_s1_allgrants) | (end_xfer_arb_share_counter_term_ram_s1 & ~ram_s1_non_bursting_master_requests);

  //ram_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ram_s1_arb_share_counter <= 0;
      else if (ram_s1_arb_counter_enable)
          ram_s1_arb_share_counter <= ram_s1_arb_share_counter_next_value;
    end


  //ram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ram_s1_slavearbiterlockenable <= 0;
      else if ((|ram_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ram_s1) | (end_xfer_arb_share_counter_term_ram_s1 & ~ram_s1_non_bursting_master_requests))
          ram_s1_slavearbiterlockenable <= |ram_s1_arb_share_counter_next_value;
    end


  //clock_crossing/m1 ram/s1 arbiterlock, which is an e_assign
  assign clock_crossing_m1_arbiterlock = ram_s1_slavearbiterlockenable & clock_crossing_m1_continuerequest;

  //ram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ram_s1_slavearbiterlockenable2 = |ram_s1_arb_share_counter_next_value;

  //clock_crossing/m1 ram/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_m1_arbiterlock2 = ram_s1_slavearbiterlockenable2 & clock_crossing_m1_continuerequest;

  //ram_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign ram_s1_any_continuerequest = 1;

  //clock_crossing_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_m1_continuerequest = 1;

  assign clock_crossing_m1_qualified_request_ram_s1 = clock_crossing_m1_requests_ram_s1 & ~((clock_crossing_m1_read & ((clock_crossing_m1_latency_counter != 0) | (1 < clock_crossing_m1_latency_counter))));
  //unique name for ram_s1_move_on_to_next_transaction, which is an e_assign
  assign ram_s1_move_on_to_next_transaction = ram_s1_readdatavalid_from_sa;

  //rdv_fifo_for_clock_crossing_m1_to_ram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_clock_crossing_m1_to_ram_s1_module rdv_fifo_for_clock_crossing_m1_to_ram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (clock_crossing_m1_granted_ram_s1),
      .data_out             (clock_crossing_m1_rdv_fifo_output_from_ram_s1),
      .empty                (),
      .fifo_contains_ones_n (clock_crossing_m1_rdv_fifo_empty_ram_s1),
      .full                 (),
      .read                 (ram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ram_s1_waits_for_read)
    );

  assign clock_crossing_m1_read_data_valid_ram_s1_shift_register = ~clock_crossing_m1_rdv_fifo_empty_ram_s1;
  //local readdatavalid clock_crossing_m1_read_data_valid_ram_s1, which is an e_mux
  assign clock_crossing_m1_read_data_valid_ram_s1 = ram_s1_readdatavalid_from_sa;

  //ram_s1_writedata mux, which is an e_mux
  assign ram_s1_writedata = clock_crossing_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_m1_granted_ram_s1 = clock_crossing_m1_qualified_request_ram_s1;

  //clock_crossing/m1 saved-grant ram/s1, which is an e_assign
  assign clock_crossing_m1_saved_grant_ram_s1 = clock_crossing_m1_requests_ram_s1;

  //allow new arb cycle for ram/s1, which is an e_assign
  assign ram_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign ram_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign ram_s1_master_qreq_vector = 1;

  //assign ram_s1_resetrequest_n_from_sa = ram_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ram_s1_resetrequest_n_from_sa = ram_s1_resetrequest_n;

  //ram_s1_firsttransfer first transaction, which is an e_assign
  assign ram_s1_firsttransfer = ram_s1_begins_xfer ? ram_s1_unreg_firsttransfer : ram_s1_reg_firsttransfer;

  //ram_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ram_s1_unreg_firsttransfer = ~(ram_s1_slavearbiterlockenable & ram_s1_any_continuerequest);

  //ram_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ram_s1_reg_firsttransfer <= 1'b1;
      else if (ram_s1_begins_xfer)
          ram_s1_reg_firsttransfer <= ram_s1_unreg_firsttransfer;
    end


  //ram_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign ram_s1_next_bbt_burstcount = ((((ram_s1_write) && (ram_s1_bbt_burstcounter == 0))))? (ram_s1_burstcount - 1) :
    ((((ram_s1_read) && (ram_s1_bbt_burstcounter == 0))))? 0 :
    (ram_s1_bbt_burstcounter - 1);

  //ram_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ram_s1_bbt_burstcounter <= 0;
      else if (ram_s1_begins_xfer)
          ram_s1_bbt_burstcounter <= ram_s1_next_bbt_burstcount;
    end


  //ram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ram_s1_beginbursttransfer_internal = ram_s1_begins_xfer & (ram_s1_bbt_burstcounter == 0);

  //ram/s1 begin burst transfer to slave, which is an e_assign
  assign ram_s1_beginbursttransfer = ram_s1_beginbursttransfer_internal;

  //ram_s1_read assignment, which is an e_mux
  assign ram_s1_read = clock_crossing_m1_granted_ram_s1 & clock_crossing_m1_read;

  //ram_s1_write assignment, which is an e_mux
  assign ram_s1_write = clock_crossing_m1_granted_ram_s1 & clock_crossing_m1_write;

  assign shifted_address_to_ram_s1_from_clock_crossing_m1 = clock_crossing_m1_address_to_slave;
  //ram_s1_address mux, which is an e_mux
  assign ram_s1_address = shifted_address_to_ram_s1_from_clock_crossing_m1 >> 2;

  //d1_ram_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ram_s1_end_xfer <= 1;
      else 
        d1_ram_s1_end_xfer <= ram_s1_end_xfer;
    end


  //ram_s1_waits_for_read in a cycle, which is an e_mux
  assign ram_s1_waits_for_read = ram_s1_in_a_read_cycle & ~ram_s1_waitrequest_n_from_sa;

  //ram_s1_in_a_read_cycle assignment, which is an e_assign
  assign ram_s1_in_a_read_cycle = clock_crossing_m1_granted_ram_s1 & clock_crossing_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ram_s1_in_a_read_cycle;

  //ram_s1_waits_for_write in a cycle, which is an e_mux
  assign ram_s1_waits_for_write = ram_s1_in_a_write_cycle & ~ram_s1_waitrequest_n_from_sa;

  //ram_s1_in_a_write_cycle assignment, which is an e_assign
  assign ram_s1_in_a_write_cycle = clock_crossing_m1_granted_ram_s1 & clock_crossing_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ram_s1_in_a_write_cycle;

  assign wait_for_ram_s1_counter = 0;
  //ram_s1_byteenable byte enable port mux, which is an e_mux
  assign ram_s1_byteenable = (clock_crossing_m1_granted_ram_s1)? clock_crossing_m1_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign ram_s1_burstcount = 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_reset_clk_125_domain_synch_module (
                                                        // inputs:
                                                         clk,
                                                         data_in,
                                                         reset_n,

                                                        // outputs:
                                                         data_out
                                                      )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module spi_0_spi_control_port_arbitrator (
                                           // inputs:
                                            Medipix_sopc_burst_10_downstream_address_to_slave,
                                            Medipix_sopc_burst_10_downstream_arbitrationshare,
                                            Medipix_sopc_burst_10_downstream_burstcount,
                                            Medipix_sopc_burst_10_downstream_latency_counter,
                                            Medipix_sopc_burst_10_downstream_nativeaddress,
                                            Medipix_sopc_burst_10_downstream_read,
                                            Medipix_sopc_burst_10_downstream_write,
                                            Medipix_sopc_burst_10_downstream_writedata,
                                            clk,
                                            reset_n,
                                            spi_0_spi_control_port_dataavailable,
                                            spi_0_spi_control_port_endofpacket,
                                            spi_0_spi_control_port_irq,
                                            spi_0_spi_control_port_readdata,
                                            spi_0_spi_control_port_readyfordata,

                                           // outputs:
                                            Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port,
                                            Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port,
                                            Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port,
                                            Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port,
                                            d1_spi_0_spi_control_port_end_xfer,
                                            spi_0_spi_control_port_address,
                                            spi_0_spi_control_port_chipselect,
                                            spi_0_spi_control_port_dataavailable_from_sa,
                                            spi_0_spi_control_port_endofpacket_from_sa,
                                            spi_0_spi_control_port_irq_from_sa,
                                            spi_0_spi_control_port_read_n,
                                            spi_0_spi_control_port_readdata_from_sa,
                                            spi_0_spi_control_port_readyfordata_from_sa,
                                            spi_0_spi_control_port_reset_n,
                                            spi_0_spi_control_port_write_n,
                                            spi_0_spi_control_port_writedata
                                         )
;

  output           Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port;
  output           Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port;
  output           Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port;
  output           Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port;
  output           d1_spi_0_spi_control_port_end_xfer;
  output  [  2: 0] spi_0_spi_control_port_address;
  output           spi_0_spi_control_port_chipselect;
  output           spi_0_spi_control_port_dataavailable_from_sa;
  output           spi_0_spi_control_port_endofpacket_from_sa;
  output           spi_0_spi_control_port_irq_from_sa;
  output           spi_0_spi_control_port_read_n;
  output  [ 15: 0] spi_0_spi_control_port_readdata_from_sa;
  output           spi_0_spi_control_port_readyfordata_from_sa;
  output           spi_0_spi_control_port_reset_n;
  output           spi_0_spi_control_port_write_n;
  output  [ 15: 0] spi_0_spi_control_port_writedata;
  input   [  3: 0] Medipix_sopc_burst_10_downstream_address_to_slave;
  input   [  4: 0] Medipix_sopc_burst_10_downstream_arbitrationshare;
  input            Medipix_sopc_burst_10_downstream_burstcount;
  input            Medipix_sopc_burst_10_downstream_latency_counter;
  input   [  3: 0] Medipix_sopc_burst_10_downstream_nativeaddress;
  input            Medipix_sopc_burst_10_downstream_read;
  input            Medipix_sopc_burst_10_downstream_write;
  input   [ 15: 0] Medipix_sopc_burst_10_downstream_writedata;
  input            clk;
  input            reset_n;
  input            spi_0_spi_control_port_dataavailable;
  input            spi_0_spi_control_port_endofpacket;
  input            spi_0_spi_control_port_irq;
  input   [ 15: 0] spi_0_spi_control_port_readdata;
  input            spi_0_spi_control_port_readyfordata;

  wire             Medipix_sopc_burst_10_downstream_arbiterlock;
  wire             Medipix_sopc_burst_10_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_10_downstream_continuerequest;
  wire             Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_saved_grant_spi_0_spi_control_port;
  reg              d1_reasons_to_wait;
  reg              d1_spi_0_spi_control_port_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_spi_0_spi_control_port;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] spi_0_spi_control_port_address;
  wire             spi_0_spi_control_port_allgrants;
  wire             spi_0_spi_control_port_allow_new_arb_cycle;
  wire             spi_0_spi_control_port_any_bursting_master_saved_grant;
  wire             spi_0_spi_control_port_any_continuerequest;
  wire             spi_0_spi_control_port_arb_counter_enable;
  reg     [  4: 0] spi_0_spi_control_port_arb_share_counter;
  wire    [  4: 0] spi_0_spi_control_port_arb_share_counter_next_value;
  wire    [  4: 0] spi_0_spi_control_port_arb_share_set_values;
  wire             spi_0_spi_control_port_beginbursttransfer_internal;
  wire             spi_0_spi_control_port_begins_xfer;
  wire             spi_0_spi_control_port_chipselect;
  wire             spi_0_spi_control_port_dataavailable_from_sa;
  wire             spi_0_spi_control_port_end_xfer;
  wire             spi_0_spi_control_port_endofpacket_from_sa;
  wire             spi_0_spi_control_port_firsttransfer;
  wire             spi_0_spi_control_port_grant_vector;
  wire             spi_0_spi_control_port_in_a_read_cycle;
  wire             spi_0_spi_control_port_in_a_write_cycle;
  wire             spi_0_spi_control_port_irq_from_sa;
  wire             spi_0_spi_control_port_master_qreq_vector;
  wire             spi_0_spi_control_port_non_bursting_master_requests;
  wire             spi_0_spi_control_port_read_n;
  wire    [ 15: 0] spi_0_spi_control_port_readdata_from_sa;
  wire             spi_0_spi_control_port_readyfordata_from_sa;
  reg              spi_0_spi_control_port_reg_firsttransfer;
  wire             spi_0_spi_control_port_reset_n;
  reg              spi_0_spi_control_port_slavearbiterlockenable;
  wire             spi_0_spi_control_port_slavearbiterlockenable2;
  wire             spi_0_spi_control_port_unreg_firsttransfer;
  wire             spi_0_spi_control_port_waits_for_read;
  wire             spi_0_spi_control_port_waits_for_write;
  wire             spi_0_spi_control_port_write_n;
  wire    [ 15: 0] spi_0_spi_control_port_writedata;
  wire             wait_for_spi_0_spi_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~spi_0_spi_control_port_end_xfer;
    end


  assign spi_0_spi_control_port_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port));
  //assign spi_0_spi_control_port_readdata_from_sa = spi_0_spi_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign spi_0_spi_control_port_readdata_from_sa = spi_0_spi_control_port_readdata;

  assign Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port = (1) & (Medipix_sopc_burst_10_downstream_read | Medipix_sopc_burst_10_downstream_write);
  //assign spi_0_spi_control_port_dataavailable_from_sa = spi_0_spi_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign spi_0_spi_control_port_dataavailable_from_sa = spi_0_spi_control_port_dataavailable;

  //assign spi_0_spi_control_port_readyfordata_from_sa = spi_0_spi_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign spi_0_spi_control_port_readyfordata_from_sa = spi_0_spi_control_port_readyfordata;

  //spi_0_spi_control_port_arb_share_counter set values, which is an e_mux
  assign spi_0_spi_control_port_arb_share_set_values = (Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port)? Medipix_sopc_burst_10_downstream_arbitrationshare :
    1;

  //spi_0_spi_control_port_non_bursting_master_requests mux, which is an e_mux
  assign spi_0_spi_control_port_non_bursting_master_requests = 0;

  //spi_0_spi_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign spi_0_spi_control_port_any_bursting_master_saved_grant = Medipix_sopc_burst_10_downstream_saved_grant_spi_0_spi_control_port;

  //spi_0_spi_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign spi_0_spi_control_port_arb_share_counter_next_value = spi_0_spi_control_port_firsttransfer ? (spi_0_spi_control_port_arb_share_set_values - 1) : |spi_0_spi_control_port_arb_share_counter ? (spi_0_spi_control_port_arb_share_counter - 1) : 0;

  //spi_0_spi_control_port_allgrants all slave grants, which is an e_mux
  assign spi_0_spi_control_port_allgrants = |spi_0_spi_control_port_grant_vector;

  //spi_0_spi_control_port_end_xfer assignment, which is an e_assign
  assign spi_0_spi_control_port_end_xfer = ~(spi_0_spi_control_port_waits_for_read | spi_0_spi_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_spi_0_spi_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_spi_0_spi_control_port = spi_0_spi_control_port_end_xfer & (~spi_0_spi_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //spi_0_spi_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign spi_0_spi_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_spi_0_spi_control_port & spi_0_spi_control_port_allgrants) | (end_xfer_arb_share_counter_term_spi_0_spi_control_port & ~spi_0_spi_control_port_non_bursting_master_requests);

  //spi_0_spi_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          spi_0_spi_control_port_arb_share_counter <= 0;
      else if (spi_0_spi_control_port_arb_counter_enable)
          spi_0_spi_control_port_arb_share_counter <= spi_0_spi_control_port_arb_share_counter_next_value;
    end


  //spi_0_spi_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          spi_0_spi_control_port_slavearbiterlockenable <= 0;
      else if ((|spi_0_spi_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_spi_0_spi_control_port) | (end_xfer_arb_share_counter_term_spi_0_spi_control_port & ~spi_0_spi_control_port_non_bursting_master_requests))
          spi_0_spi_control_port_slavearbiterlockenable <= |spi_0_spi_control_port_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_10/downstream spi_0/spi_control_port arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_arbiterlock = spi_0_spi_control_port_slavearbiterlockenable & Medipix_sopc_burst_10_downstream_continuerequest;

  //spi_0_spi_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign spi_0_spi_control_port_slavearbiterlockenable2 = |spi_0_spi_control_port_arb_share_counter_next_value;

  //Medipix_sopc_burst_10/downstream spi_0/spi_control_port arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_arbiterlock2 = spi_0_spi_control_port_slavearbiterlockenable2 & Medipix_sopc_burst_10_downstream_continuerequest;

  //spi_0_spi_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  assign spi_0_spi_control_port_any_continuerequest = 1;

  //Medipix_sopc_burst_10_downstream_continuerequest continued request, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_continuerequest = 1;

  assign Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port = Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port & ~((Medipix_sopc_burst_10_downstream_read & ((Medipix_sopc_burst_10_downstream_latency_counter != 0))));
  //local readdatavalid Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port, which is an e_mux
  assign Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port = Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port & Medipix_sopc_burst_10_downstream_read & ~spi_0_spi_control_port_waits_for_read;

  //spi_0_spi_control_port_writedata mux, which is an e_mux
  assign spi_0_spi_control_port_writedata = Medipix_sopc_burst_10_downstream_writedata;

  //assign spi_0_spi_control_port_endofpacket_from_sa = spi_0_spi_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign spi_0_spi_control_port_endofpacket_from_sa = spi_0_spi_control_port_endofpacket;

  //master is always granted when requested
  assign Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port = Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port;

  //Medipix_sopc_burst_10/downstream saved-grant spi_0/spi_control_port, which is an e_assign
  assign Medipix_sopc_burst_10_downstream_saved_grant_spi_0_spi_control_port = Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port;

  //allow new arb cycle for spi_0/spi_control_port, which is an e_assign
  assign spi_0_spi_control_port_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign spi_0_spi_control_port_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign spi_0_spi_control_port_master_qreq_vector = 1;

  //spi_0_spi_control_port_reset_n assignment, which is an e_assign
  assign spi_0_spi_control_port_reset_n = reset_n;

  assign spi_0_spi_control_port_chipselect = Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port;
  //spi_0_spi_control_port_firsttransfer first transaction, which is an e_assign
  assign spi_0_spi_control_port_firsttransfer = spi_0_spi_control_port_begins_xfer ? spi_0_spi_control_port_unreg_firsttransfer : spi_0_spi_control_port_reg_firsttransfer;

  //spi_0_spi_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign spi_0_spi_control_port_unreg_firsttransfer = ~(spi_0_spi_control_port_slavearbiterlockenable & spi_0_spi_control_port_any_continuerequest);

  //spi_0_spi_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          spi_0_spi_control_port_reg_firsttransfer <= 1'b1;
      else if (spi_0_spi_control_port_begins_xfer)
          spi_0_spi_control_port_reg_firsttransfer <= spi_0_spi_control_port_unreg_firsttransfer;
    end


  //spi_0_spi_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign spi_0_spi_control_port_beginbursttransfer_internal = spi_0_spi_control_port_begins_xfer;

  //~spi_0_spi_control_port_read_n assignment, which is an e_mux
  assign spi_0_spi_control_port_read_n = ~(Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port & Medipix_sopc_burst_10_downstream_read);

  //~spi_0_spi_control_port_write_n assignment, which is an e_mux
  assign spi_0_spi_control_port_write_n = ~(Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port & Medipix_sopc_burst_10_downstream_write);

  //spi_0_spi_control_port_address mux, which is an e_mux
  assign spi_0_spi_control_port_address = Medipix_sopc_burst_10_downstream_nativeaddress;

  //d1_spi_0_spi_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_spi_0_spi_control_port_end_xfer <= 1;
      else 
        d1_spi_0_spi_control_port_end_xfer <= spi_0_spi_control_port_end_xfer;
    end


  //spi_0_spi_control_port_waits_for_read in a cycle, which is an e_mux
  assign spi_0_spi_control_port_waits_for_read = spi_0_spi_control_port_in_a_read_cycle & spi_0_spi_control_port_begins_xfer;

  //spi_0_spi_control_port_in_a_read_cycle assignment, which is an e_assign
  assign spi_0_spi_control_port_in_a_read_cycle = Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port & Medipix_sopc_burst_10_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = spi_0_spi_control_port_in_a_read_cycle;

  //spi_0_spi_control_port_waits_for_write in a cycle, which is an e_mux
  assign spi_0_spi_control_port_waits_for_write = spi_0_spi_control_port_in_a_write_cycle & spi_0_spi_control_port_begins_xfer;

  //spi_0_spi_control_port_in_a_write_cycle assignment, which is an e_assign
  assign spi_0_spi_control_port_in_a_write_cycle = Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port & Medipix_sopc_burst_10_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = spi_0_spi_control_port_in_a_write_cycle;

  assign wait_for_spi_0_spi_control_port_counter = 0;
  //assign spi_0_spi_control_port_irq_from_sa = spi_0_spi_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign spi_0_spi_control_port_irq_from_sa = spi_0_spi_control_port_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //spi_0/spi_control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_10/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port && (Medipix_sopc_burst_10_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_10/downstream drove 0 on its 'arbitrationshare' port while accessing slave spi_0/spi_control_port", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_10/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port && (Medipix_sopc_burst_10_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_10/downstream drove 0 on its 'burstcount' port while accessing slave spi_0/spi_control_port", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sys_clk_freq_s1_arbitrator (
                                    // inputs:
                                     Medipix_sopc_burst_3_downstream_address_to_slave,
                                     Medipix_sopc_burst_3_downstream_arbitrationshare,
                                     Medipix_sopc_burst_3_downstream_burstcount,
                                     Medipix_sopc_burst_3_downstream_latency_counter,
                                     Medipix_sopc_burst_3_downstream_nativeaddress,
                                     Medipix_sopc_burst_3_downstream_read,
                                     Medipix_sopc_burst_3_downstream_write,
                                     Medipix_sopc_burst_3_downstream_writedata,
                                     clk,
                                     reset_n,
                                     sys_clk_freq_s1_irq,
                                     sys_clk_freq_s1_readdata,

                                    // outputs:
                                     Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1,
                                     Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1,
                                     Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1,
                                     Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1,
                                     d1_sys_clk_freq_s1_end_xfer,
                                     sys_clk_freq_s1_address,
                                     sys_clk_freq_s1_chipselect,
                                     sys_clk_freq_s1_irq_from_sa,
                                     sys_clk_freq_s1_readdata_from_sa,
                                     sys_clk_freq_s1_reset_n,
                                     sys_clk_freq_s1_write_n,
                                     sys_clk_freq_s1_writedata
                                  )
;

  output           Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1;
  output           Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1;
  output           Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1;
  output           Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1;
  output           d1_sys_clk_freq_s1_end_xfer;
  output  [  2: 0] sys_clk_freq_s1_address;
  output           sys_clk_freq_s1_chipselect;
  output           sys_clk_freq_s1_irq_from_sa;
  output  [ 15: 0] sys_clk_freq_s1_readdata_from_sa;
  output           sys_clk_freq_s1_reset_n;
  output           sys_clk_freq_s1_write_n;
  output  [ 15: 0] sys_clk_freq_s1_writedata;
  input   [  3: 0] Medipix_sopc_burst_3_downstream_address_to_slave;
  input   [  4: 0] Medipix_sopc_burst_3_downstream_arbitrationshare;
  input            Medipix_sopc_burst_3_downstream_burstcount;
  input            Medipix_sopc_burst_3_downstream_latency_counter;
  input   [  3: 0] Medipix_sopc_burst_3_downstream_nativeaddress;
  input            Medipix_sopc_burst_3_downstream_read;
  input            Medipix_sopc_burst_3_downstream_write;
  input   [ 15: 0] Medipix_sopc_burst_3_downstream_writedata;
  input            clk;
  input            reset_n;
  input            sys_clk_freq_s1_irq;
  input   [ 15: 0] sys_clk_freq_s1_readdata;

  wire             Medipix_sopc_burst_3_downstream_arbiterlock;
  wire             Medipix_sopc_burst_3_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_3_downstream_continuerequest;
  wire             Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_saved_grant_sys_clk_freq_s1;
  reg              d1_reasons_to_wait;
  reg              d1_sys_clk_freq_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sys_clk_freq_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] sys_clk_freq_s1_address;
  wire             sys_clk_freq_s1_allgrants;
  wire             sys_clk_freq_s1_allow_new_arb_cycle;
  wire             sys_clk_freq_s1_any_bursting_master_saved_grant;
  wire             sys_clk_freq_s1_any_continuerequest;
  wire             sys_clk_freq_s1_arb_counter_enable;
  reg     [  4: 0] sys_clk_freq_s1_arb_share_counter;
  wire    [  4: 0] sys_clk_freq_s1_arb_share_counter_next_value;
  wire    [  4: 0] sys_clk_freq_s1_arb_share_set_values;
  wire             sys_clk_freq_s1_beginbursttransfer_internal;
  wire             sys_clk_freq_s1_begins_xfer;
  wire             sys_clk_freq_s1_chipselect;
  wire             sys_clk_freq_s1_end_xfer;
  wire             sys_clk_freq_s1_firsttransfer;
  wire             sys_clk_freq_s1_grant_vector;
  wire             sys_clk_freq_s1_in_a_read_cycle;
  wire             sys_clk_freq_s1_in_a_write_cycle;
  wire             sys_clk_freq_s1_irq_from_sa;
  wire             sys_clk_freq_s1_master_qreq_vector;
  wire             sys_clk_freq_s1_non_bursting_master_requests;
  wire    [ 15: 0] sys_clk_freq_s1_readdata_from_sa;
  reg              sys_clk_freq_s1_reg_firsttransfer;
  wire             sys_clk_freq_s1_reset_n;
  reg              sys_clk_freq_s1_slavearbiterlockenable;
  wire             sys_clk_freq_s1_slavearbiterlockenable2;
  wire             sys_clk_freq_s1_unreg_firsttransfer;
  wire             sys_clk_freq_s1_waits_for_read;
  wire             sys_clk_freq_s1_waits_for_write;
  wire             sys_clk_freq_s1_write_n;
  wire    [ 15: 0] sys_clk_freq_s1_writedata;
  wire             wait_for_sys_clk_freq_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sys_clk_freq_s1_end_xfer;
    end


  assign sys_clk_freq_s1_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1));
  //assign sys_clk_freq_s1_readdata_from_sa = sys_clk_freq_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_clk_freq_s1_readdata_from_sa = sys_clk_freq_s1_readdata;

  assign Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1 = (1) & (Medipix_sopc_burst_3_downstream_read | Medipix_sopc_burst_3_downstream_write);
  //sys_clk_freq_s1_arb_share_counter set values, which is an e_mux
  assign sys_clk_freq_s1_arb_share_set_values = (Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1)? Medipix_sopc_burst_3_downstream_arbitrationshare :
    1;

  //sys_clk_freq_s1_non_bursting_master_requests mux, which is an e_mux
  assign sys_clk_freq_s1_non_bursting_master_requests = 0;

  //sys_clk_freq_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sys_clk_freq_s1_any_bursting_master_saved_grant = Medipix_sopc_burst_3_downstream_saved_grant_sys_clk_freq_s1;

  //sys_clk_freq_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sys_clk_freq_s1_arb_share_counter_next_value = sys_clk_freq_s1_firsttransfer ? (sys_clk_freq_s1_arb_share_set_values - 1) : |sys_clk_freq_s1_arb_share_counter ? (sys_clk_freq_s1_arb_share_counter - 1) : 0;

  //sys_clk_freq_s1_allgrants all slave grants, which is an e_mux
  assign sys_clk_freq_s1_allgrants = |sys_clk_freq_s1_grant_vector;

  //sys_clk_freq_s1_end_xfer assignment, which is an e_assign
  assign sys_clk_freq_s1_end_xfer = ~(sys_clk_freq_s1_waits_for_read | sys_clk_freq_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sys_clk_freq_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sys_clk_freq_s1 = sys_clk_freq_s1_end_xfer & (~sys_clk_freq_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sys_clk_freq_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sys_clk_freq_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sys_clk_freq_s1 & sys_clk_freq_s1_allgrants) | (end_xfer_arb_share_counter_term_sys_clk_freq_s1 & ~sys_clk_freq_s1_non_bursting_master_requests);

  //sys_clk_freq_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_freq_s1_arb_share_counter <= 0;
      else if (sys_clk_freq_s1_arb_counter_enable)
          sys_clk_freq_s1_arb_share_counter <= sys_clk_freq_s1_arb_share_counter_next_value;
    end


  //sys_clk_freq_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_freq_s1_slavearbiterlockenable <= 0;
      else if ((|sys_clk_freq_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sys_clk_freq_s1) | (end_xfer_arb_share_counter_term_sys_clk_freq_s1 & ~sys_clk_freq_s1_non_bursting_master_requests))
          sys_clk_freq_s1_slavearbiterlockenable <= |sys_clk_freq_s1_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_3/downstream sys_clk_freq/s1 arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_arbiterlock = sys_clk_freq_s1_slavearbiterlockenable & Medipix_sopc_burst_3_downstream_continuerequest;

  //sys_clk_freq_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sys_clk_freq_s1_slavearbiterlockenable2 = |sys_clk_freq_s1_arb_share_counter_next_value;

  //Medipix_sopc_burst_3/downstream sys_clk_freq/s1 arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_arbiterlock2 = sys_clk_freq_s1_slavearbiterlockenable2 & Medipix_sopc_burst_3_downstream_continuerequest;

  //sys_clk_freq_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sys_clk_freq_s1_any_continuerequest = 1;

  //Medipix_sopc_burst_3_downstream_continuerequest continued request, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_continuerequest = 1;

  assign Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1 = Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1 & ~((Medipix_sopc_burst_3_downstream_read & ((Medipix_sopc_burst_3_downstream_latency_counter != 0))));
  //local readdatavalid Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1, which is an e_mux
  assign Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1 = Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1 & Medipix_sopc_burst_3_downstream_read & ~sys_clk_freq_s1_waits_for_read;

  //sys_clk_freq_s1_writedata mux, which is an e_mux
  assign sys_clk_freq_s1_writedata = Medipix_sopc_burst_3_downstream_writedata;

  //master is always granted when requested
  assign Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1 = Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1;

  //Medipix_sopc_burst_3/downstream saved-grant sys_clk_freq/s1, which is an e_assign
  assign Medipix_sopc_burst_3_downstream_saved_grant_sys_clk_freq_s1 = Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1;

  //allow new arb cycle for sys_clk_freq/s1, which is an e_assign
  assign sys_clk_freq_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sys_clk_freq_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sys_clk_freq_s1_master_qreq_vector = 1;

  //sys_clk_freq_s1_reset_n assignment, which is an e_assign
  assign sys_clk_freq_s1_reset_n = reset_n;

  assign sys_clk_freq_s1_chipselect = Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1;
  //sys_clk_freq_s1_firsttransfer first transaction, which is an e_assign
  assign sys_clk_freq_s1_firsttransfer = sys_clk_freq_s1_begins_xfer ? sys_clk_freq_s1_unreg_firsttransfer : sys_clk_freq_s1_reg_firsttransfer;

  //sys_clk_freq_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sys_clk_freq_s1_unreg_firsttransfer = ~(sys_clk_freq_s1_slavearbiterlockenable & sys_clk_freq_s1_any_continuerequest);

  //sys_clk_freq_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_freq_s1_reg_firsttransfer <= 1'b1;
      else if (sys_clk_freq_s1_begins_xfer)
          sys_clk_freq_s1_reg_firsttransfer <= sys_clk_freq_s1_unreg_firsttransfer;
    end


  //sys_clk_freq_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sys_clk_freq_s1_beginbursttransfer_internal = sys_clk_freq_s1_begins_xfer;

  //~sys_clk_freq_s1_write_n assignment, which is an e_mux
  assign sys_clk_freq_s1_write_n = ~(Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1 & Medipix_sopc_burst_3_downstream_write);

  //sys_clk_freq_s1_address mux, which is an e_mux
  assign sys_clk_freq_s1_address = Medipix_sopc_burst_3_downstream_nativeaddress;

  //d1_sys_clk_freq_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sys_clk_freq_s1_end_xfer <= 1;
      else 
        d1_sys_clk_freq_s1_end_xfer <= sys_clk_freq_s1_end_xfer;
    end


  //sys_clk_freq_s1_waits_for_read in a cycle, which is an e_mux
  assign sys_clk_freq_s1_waits_for_read = sys_clk_freq_s1_in_a_read_cycle & sys_clk_freq_s1_begins_xfer;

  //sys_clk_freq_s1_in_a_read_cycle assignment, which is an e_assign
  assign sys_clk_freq_s1_in_a_read_cycle = Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1 & Medipix_sopc_burst_3_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sys_clk_freq_s1_in_a_read_cycle;

  //sys_clk_freq_s1_waits_for_write in a cycle, which is an e_mux
  assign sys_clk_freq_s1_waits_for_write = sys_clk_freq_s1_in_a_write_cycle & 0;

  //sys_clk_freq_s1_in_a_write_cycle assignment, which is an e_assign
  assign sys_clk_freq_s1_in_a_write_cycle = Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1 & Medipix_sopc_burst_3_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sys_clk_freq_s1_in_a_write_cycle;

  assign wait_for_sys_clk_freq_s1_counter = 0;
  //assign sys_clk_freq_s1_irq_from_sa = sys_clk_freq_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_clk_freq_s1_irq_from_sa = sys_clk_freq_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sys_clk_freq/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_3/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1 && (Medipix_sopc_burst_3_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_3/downstream drove 0 on its 'arbitrationshare' port while accessing slave sys_clk_freq/s1", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_3/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1 && (Medipix_sopc_burst_3_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_3/downstream drove 0 on its 'burstcount' port while accessing slave sys_clk_freq/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tx_table_avalon_slave_0_arbitrator (
                                            // inputs:
                                             Medipix_sopc_burst_9_downstream_address_to_slave,
                                             Medipix_sopc_burst_9_downstream_arbitrationshare,
                                             Medipix_sopc_burst_9_downstream_burstcount,
                                             Medipix_sopc_burst_9_downstream_latency_counter,
                                             Medipix_sopc_burst_9_downstream_read,
                                             Medipix_sopc_burst_9_downstream_write,
                                             Medipix_sopc_burst_9_downstream_writedata,
                                             clk,
                                             reset_n,
                                             tx_table_avalon_slave_0_readdata,

                                            // outputs:
                                             Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0,
                                             Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0,
                                             Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0,
                                             Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0,
                                             d1_tx_table_avalon_slave_0_end_xfer,
                                             tx_table_avalon_slave_0_address,
                                             tx_table_avalon_slave_0_chipselect,
                                             tx_table_avalon_slave_0_read,
                                             tx_table_avalon_slave_0_readdata_from_sa,
                                             tx_table_avalon_slave_0_reset_n,
                                             tx_table_avalon_slave_0_write,
                                             tx_table_avalon_slave_0_writedata
                                          )
;

  output           Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0;
  output           Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0;
  output           Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0;
  output           Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0;
  output           d1_tx_table_avalon_slave_0_end_xfer;
  output  [  1: 0] tx_table_avalon_slave_0_address;
  output           tx_table_avalon_slave_0_chipselect;
  output           tx_table_avalon_slave_0_read;
  output  [ 31: 0] tx_table_avalon_slave_0_readdata_from_sa;
  output           tx_table_avalon_slave_0_reset_n;
  output           tx_table_avalon_slave_0_write;
  output  [ 31: 0] tx_table_avalon_slave_0_writedata;
  input   [  3: 0] Medipix_sopc_burst_9_downstream_address_to_slave;
  input   [  3: 0] Medipix_sopc_burst_9_downstream_arbitrationshare;
  input            Medipix_sopc_burst_9_downstream_burstcount;
  input            Medipix_sopc_burst_9_downstream_latency_counter;
  input            Medipix_sopc_burst_9_downstream_read;
  input            Medipix_sopc_burst_9_downstream_write;
  input   [ 31: 0] Medipix_sopc_burst_9_downstream_writedata;
  input            clk;
  input            reset_n;
  input   [ 31: 0] tx_table_avalon_slave_0_readdata;

  wire             Medipix_sopc_burst_9_downstream_arbiterlock;
  wire             Medipix_sopc_burst_9_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_9_downstream_continuerequest;
  wire             Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_saved_grant_tx_table_avalon_slave_0;
  reg              d1_reasons_to_wait;
  reg              d1_tx_table_avalon_slave_0_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tx_table_avalon_slave_0;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  3: 0] shifted_address_to_tx_table_avalon_slave_0_from_Medipix_sopc_burst_9_downstream;
  wire    [  1: 0] tx_table_avalon_slave_0_address;
  wire             tx_table_avalon_slave_0_allgrants;
  wire             tx_table_avalon_slave_0_allow_new_arb_cycle;
  wire             tx_table_avalon_slave_0_any_bursting_master_saved_grant;
  wire             tx_table_avalon_slave_0_any_continuerequest;
  wire             tx_table_avalon_slave_0_arb_counter_enable;
  reg     [  3: 0] tx_table_avalon_slave_0_arb_share_counter;
  wire    [  3: 0] tx_table_avalon_slave_0_arb_share_counter_next_value;
  wire    [  3: 0] tx_table_avalon_slave_0_arb_share_set_values;
  wire             tx_table_avalon_slave_0_beginbursttransfer_internal;
  wire             tx_table_avalon_slave_0_begins_xfer;
  wire             tx_table_avalon_slave_0_chipselect;
  wire             tx_table_avalon_slave_0_end_xfer;
  wire             tx_table_avalon_slave_0_firsttransfer;
  wire             tx_table_avalon_slave_0_grant_vector;
  wire             tx_table_avalon_slave_0_in_a_read_cycle;
  wire             tx_table_avalon_slave_0_in_a_write_cycle;
  wire             tx_table_avalon_slave_0_master_qreq_vector;
  wire             tx_table_avalon_slave_0_non_bursting_master_requests;
  wire             tx_table_avalon_slave_0_read;
  wire    [ 31: 0] tx_table_avalon_slave_0_readdata_from_sa;
  reg              tx_table_avalon_slave_0_reg_firsttransfer;
  wire             tx_table_avalon_slave_0_reset_n;
  reg              tx_table_avalon_slave_0_slavearbiterlockenable;
  wire             tx_table_avalon_slave_0_slavearbiterlockenable2;
  wire             tx_table_avalon_slave_0_unreg_firsttransfer;
  wire             tx_table_avalon_slave_0_waits_for_read;
  wire             tx_table_avalon_slave_0_waits_for_write;
  wire             tx_table_avalon_slave_0_write;
  wire    [ 31: 0] tx_table_avalon_slave_0_writedata;
  wire             wait_for_tx_table_avalon_slave_0_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tx_table_avalon_slave_0_end_xfer;
    end


  assign tx_table_avalon_slave_0_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0));
  //assign tx_table_avalon_slave_0_readdata_from_sa = tx_table_avalon_slave_0_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tx_table_avalon_slave_0_readdata_from_sa = tx_table_avalon_slave_0_readdata;

  assign Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0 = (1) & (Medipix_sopc_burst_9_downstream_read | Medipix_sopc_burst_9_downstream_write);
  //tx_table_avalon_slave_0_arb_share_counter set values, which is an e_mux
  assign tx_table_avalon_slave_0_arb_share_set_values = (Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0)? Medipix_sopc_burst_9_downstream_arbitrationshare :
    1;

  //tx_table_avalon_slave_0_non_bursting_master_requests mux, which is an e_mux
  assign tx_table_avalon_slave_0_non_bursting_master_requests = 0;

  //tx_table_avalon_slave_0_any_bursting_master_saved_grant mux, which is an e_mux
  assign tx_table_avalon_slave_0_any_bursting_master_saved_grant = Medipix_sopc_burst_9_downstream_saved_grant_tx_table_avalon_slave_0;

  //tx_table_avalon_slave_0_arb_share_counter_next_value assignment, which is an e_assign
  assign tx_table_avalon_slave_0_arb_share_counter_next_value = tx_table_avalon_slave_0_firsttransfer ? (tx_table_avalon_slave_0_arb_share_set_values - 1) : |tx_table_avalon_slave_0_arb_share_counter ? (tx_table_avalon_slave_0_arb_share_counter - 1) : 0;

  //tx_table_avalon_slave_0_allgrants all slave grants, which is an e_mux
  assign tx_table_avalon_slave_0_allgrants = |tx_table_avalon_slave_0_grant_vector;

  //tx_table_avalon_slave_0_end_xfer assignment, which is an e_assign
  assign tx_table_avalon_slave_0_end_xfer = ~(tx_table_avalon_slave_0_waits_for_read | tx_table_avalon_slave_0_waits_for_write);

  //end_xfer_arb_share_counter_term_tx_table_avalon_slave_0 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tx_table_avalon_slave_0 = tx_table_avalon_slave_0_end_xfer & (~tx_table_avalon_slave_0_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tx_table_avalon_slave_0_arb_share_counter arbitration counter enable, which is an e_assign
  assign tx_table_avalon_slave_0_arb_counter_enable = (end_xfer_arb_share_counter_term_tx_table_avalon_slave_0 & tx_table_avalon_slave_0_allgrants) | (end_xfer_arb_share_counter_term_tx_table_avalon_slave_0 & ~tx_table_avalon_slave_0_non_bursting_master_requests);

  //tx_table_avalon_slave_0_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tx_table_avalon_slave_0_arb_share_counter <= 0;
      else if (tx_table_avalon_slave_0_arb_counter_enable)
          tx_table_avalon_slave_0_arb_share_counter <= tx_table_avalon_slave_0_arb_share_counter_next_value;
    end


  //tx_table_avalon_slave_0_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tx_table_avalon_slave_0_slavearbiterlockenable <= 0;
      else if ((|tx_table_avalon_slave_0_master_qreq_vector & end_xfer_arb_share_counter_term_tx_table_avalon_slave_0) | (end_xfer_arb_share_counter_term_tx_table_avalon_slave_0 & ~tx_table_avalon_slave_0_non_bursting_master_requests))
          tx_table_avalon_slave_0_slavearbiterlockenable <= |tx_table_avalon_slave_0_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_9/downstream tx_table/avalon_slave_0 arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_arbiterlock = tx_table_avalon_slave_0_slavearbiterlockenable & Medipix_sopc_burst_9_downstream_continuerequest;

  //tx_table_avalon_slave_0_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tx_table_avalon_slave_0_slavearbiterlockenable2 = |tx_table_avalon_slave_0_arb_share_counter_next_value;

  //Medipix_sopc_burst_9/downstream tx_table/avalon_slave_0 arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_arbiterlock2 = tx_table_avalon_slave_0_slavearbiterlockenable2 & Medipix_sopc_burst_9_downstream_continuerequest;

  //tx_table_avalon_slave_0_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tx_table_avalon_slave_0_any_continuerequest = 1;

  //Medipix_sopc_burst_9_downstream_continuerequest continued request, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_continuerequest = 1;

  assign Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0 = Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0 & ~((Medipix_sopc_burst_9_downstream_read & ((Medipix_sopc_burst_9_downstream_latency_counter != 0))));
  //local readdatavalid Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0, which is an e_mux
  assign Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0 = Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0 & Medipix_sopc_burst_9_downstream_read & ~tx_table_avalon_slave_0_waits_for_read;

  //tx_table_avalon_slave_0_writedata mux, which is an e_mux
  assign tx_table_avalon_slave_0_writedata = Medipix_sopc_burst_9_downstream_writedata;

  //master is always granted when requested
  assign Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0 = Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0;

  //Medipix_sopc_burst_9/downstream saved-grant tx_table/avalon_slave_0, which is an e_assign
  assign Medipix_sopc_burst_9_downstream_saved_grant_tx_table_avalon_slave_0 = Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0;

  //allow new arb cycle for tx_table/avalon_slave_0, which is an e_assign
  assign tx_table_avalon_slave_0_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tx_table_avalon_slave_0_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tx_table_avalon_slave_0_master_qreq_vector = 1;

  //tx_table_avalon_slave_0_reset_n assignment, which is an e_assign
  assign tx_table_avalon_slave_0_reset_n = reset_n;

  assign tx_table_avalon_slave_0_chipselect = Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0;
  //tx_table_avalon_slave_0_firsttransfer first transaction, which is an e_assign
  assign tx_table_avalon_slave_0_firsttransfer = tx_table_avalon_slave_0_begins_xfer ? tx_table_avalon_slave_0_unreg_firsttransfer : tx_table_avalon_slave_0_reg_firsttransfer;

  //tx_table_avalon_slave_0_unreg_firsttransfer first transaction, which is an e_assign
  assign tx_table_avalon_slave_0_unreg_firsttransfer = ~(tx_table_avalon_slave_0_slavearbiterlockenable & tx_table_avalon_slave_0_any_continuerequest);

  //tx_table_avalon_slave_0_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tx_table_avalon_slave_0_reg_firsttransfer <= 1'b1;
      else if (tx_table_avalon_slave_0_begins_xfer)
          tx_table_avalon_slave_0_reg_firsttransfer <= tx_table_avalon_slave_0_unreg_firsttransfer;
    end


  //tx_table_avalon_slave_0_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tx_table_avalon_slave_0_beginbursttransfer_internal = tx_table_avalon_slave_0_begins_xfer;

  //tx_table_avalon_slave_0_read assignment, which is an e_mux
  assign tx_table_avalon_slave_0_read = Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0 & Medipix_sopc_burst_9_downstream_read;

  //tx_table_avalon_slave_0_write assignment, which is an e_mux
  assign tx_table_avalon_slave_0_write = Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0 & Medipix_sopc_burst_9_downstream_write;

  assign shifted_address_to_tx_table_avalon_slave_0_from_Medipix_sopc_burst_9_downstream = Medipix_sopc_burst_9_downstream_address_to_slave;
  //tx_table_avalon_slave_0_address mux, which is an e_mux
  assign tx_table_avalon_slave_0_address = shifted_address_to_tx_table_avalon_slave_0_from_Medipix_sopc_burst_9_downstream >> 2;

  //d1_tx_table_avalon_slave_0_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tx_table_avalon_slave_0_end_xfer <= 1;
      else 
        d1_tx_table_avalon_slave_0_end_xfer <= tx_table_avalon_slave_0_end_xfer;
    end


  //tx_table_avalon_slave_0_waits_for_read in a cycle, which is an e_mux
  assign tx_table_avalon_slave_0_waits_for_read = tx_table_avalon_slave_0_in_a_read_cycle & tx_table_avalon_slave_0_begins_xfer;

  //tx_table_avalon_slave_0_in_a_read_cycle assignment, which is an e_assign
  assign tx_table_avalon_slave_0_in_a_read_cycle = Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0 & Medipix_sopc_burst_9_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tx_table_avalon_slave_0_in_a_read_cycle;

  //tx_table_avalon_slave_0_waits_for_write in a cycle, which is an e_mux
  assign tx_table_avalon_slave_0_waits_for_write = tx_table_avalon_slave_0_in_a_write_cycle & 0;

  //tx_table_avalon_slave_0_in_a_write_cycle assignment, which is an e_assign
  assign tx_table_avalon_slave_0_in_a_write_cycle = Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0 & Medipix_sopc_burst_9_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tx_table_avalon_slave_0_in_a_write_cycle;

  assign wait_for_tx_table_avalon_slave_0_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tx_table/avalon_slave_0 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_9/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0 && (Medipix_sopc_burst_9_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_9/downstream drove 0 on its 'arbitrationshare' port while accessing slave tx_table/avalon_slave_0", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_9/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0 && (Medipix_sopc_burst_9_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_9/downstream drove 0 on its 'burstcount' port while accessing slave tx_table/avalon_slave_0", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module uart_0_s1_arbitrator (
                              // inputs:
                               Medipix_sopc_burst_11_downstream_address_to_slave,
                               Medipix_sopc_burst_11_downstream_arbitrationshare,
                               Medipix_sopc_burst_11_downstream_burstcount,
                               Medipix_sopc_burst_11_downstream_latency_counter,
                               Medipix_sopc_burst_11_downstream_nativeaddress,
                               Medipix_sopc_burst_11_downstream_read,
                               Medipix_sopc_burst_11_downstream_write,
                               Medipix_sopc_burst_11_downstream_writedata,
                               clk,
                               reset_n,
                               uart_0_s1_dataavailable,
                               uart_0_s1_irq,
                               uart_0_s1_readdata,
                               uart_0_s1_readyfordata,

                              // outputs:
                               Medipix_sopc_burst_11_downstream_granted_uart_0_s1,
                               Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1,
                               Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1,
                               Medipix_sopc_burst_11_downstream_requests_uart_0_s1,
                               d1_uart_0_s1_end_xfer,
                               uart_0_s1_address,
                               uart_0_s1_begintransfer,
                               uart_0_s1_chipselect,
                               uart_0_s1_dataavailable_from_sa,
                               uart_0_s1_irq_from_sa,
                               uart_0_s1_read_n,
                               uart_0_s1_readdata_from_sa,
                               uart_0_s1_readyfordata_from_sa,
                               uart_0_s1_reset_n,
                               uart_0_s1_write_n,
                               uart_0_s1_writedata
                            )
;

  output           Medipix_sopc_burst_11_downstream_granted_uart_0_s1;
  output           Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1;
  output           Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1;
  output           Medipix_sopc_burst_11_downstream_requests_uart_0_s1;
  output           d1_uart_0_s1_end_xfer;
  output  [  2: 0] uart_0_s1_address;
  output           uart_0_s1_begintransfer;
  output           uart_0_s1_chipselect;
  output           uart_0_s1_dataavailable_from_sa;
  output           uart_0_s1_irq_from_sa;
  output           uart_0_s1_read_n;
  output  [ 15: 0] uart_0_s1_readdata_from_sa;
  output           uart_0_s1_readyfordata_from_sa;
  output           uart_0_s1_reset_n;
  output           uart_0_s1_write_n;
  output  [ 15: 0] uart_0_s1_writedata;
  input   [  3: 0] Medipix_sopc_burst_11_downstream_address_to_slave;
  input   [  4: 0] Medipix_sopc_burst_11_downstream_arbitrationshare;
  input            Medipix_sopc_burst_11_downstream_burstcount;
  input            Medipix_sopc_burst_11_downstream_latency_counter;
  input   [  3: 0] Medipix_sopc_burst_11_downstream_nativeaddress;
  input            Medipix_sopc_burst_11_downstream_read;
  input            Medipix_sopc_burst_11_downstream_write;
  input   [ 15: 0] Medipix_sopc_burst_11_downstream_writedata;
  input            clk;
  input            reset_n;
  input            uart_0_s1_dataavailable;
  input            uart_0_s1_irq;
  input   [ 15: 0] uart_0_s1_readdata;
  input            uart_0_s1_readyfordata;

  wire             Medipix_sopc_burst_11_downstream_arbiterlock;
  wire             Medipix_sopc_burst_11_downstream_arbiterlock2;
  wire             Medipix_sopc_burst_11_downstream_continuerequest;
  wire             Medipix_sopc_burst_11_downstream_granted_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_requests_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_saved_grant_uart_0_s1;
  reg              d1_reasons_to_wait;
  reg              d1_uart_0_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_uart_0_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] uart_0_s1_address;
  wire             uart_0_s1_allgrants;
  wire             uart_0_s1_allow_new_arb_cycle;
  wire             uart_0_s1_any_bursting_master_saved_grant;
  wire             uart_0_s1_any_continuerequest;
  wire             uart_0_s1_arb_counter_enable;
  reg     [  4: 0] uart_0_s1_arb_share_counter;
  wire    [  4: 0] uart_0_s1_arb_share_counter_next_value;
  wire    [  4: 0] uart_0_s1_arb_share_set_values;
  wire             uart_0_s1_beginbursttransfer_internal;
  wire             uart_0_s1_begins_xfer;
  wire             uart_0_s1_begintransfer;
  wire             uart_0_s1_chipselect;
  wire             uart_0_s1_dataavailable_from_sa;
  wire             uart_0_s1_end_xfer;
  wire             uart_0_s1_firsttransfer;
  wire             uart_0_s1_grant_vector;
  wire             uart_0_s1_in_a_read_cycle;
  wire             uart_0_s1_in_a_write_cycle;
  wire             uart_0_s1_irq_from_sa;
  wire             uart_0_s1_master_qreq_vector;
  wire             uart_0_s1_non_bursting_master_requests;
  wire             uart_0_s1_read_n;
  wire    [ 15: 0] uart_0_s1_readdata_from_sa;
  wire             uart_0_s1_readyfordata_from_sa;
  reg              uart_0_s1_reg_firsttransfer;
  wire             uart_0_s1_reset_n;
  reg              uart_0_s1_slavearbiterlockenable;
  wire             uart_0_s1_slavearbiterlockenable2;
  wire             uart_0_s1_unreg_firsttransfer;
  wire             uart_0_s1_waits_for_read;
  wire             uart_0_s1_waits_for_write;
  wire             uart_0_s1_write_n;
  wire    [ 15: 0] uart_0_s1_writedata;
  wire             wait_for_uart_0_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~uart_0_s1_end_xfer;
    end


  assign uart_0_s1_begins_xfer = ~d1_reasons_to_wait & ((Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1));
  //assign uart_0_s1_readdata_from_sa = uart_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_0_s1_readdata_from_sa = uart_0_s1_readdata;

  assign Medipix_sopc_burst_11_downstream_requests_uart_0_s1 = (1) & (Medipix_sopc_burst_11_downstream_read | Medipix_sopc_burst_11_downstream_write);
  //assign uart_0_s1_dataavailable_from_sa = uart_0_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_0_s1_dataavailable_from_sa = uart_0_s1_dataavailable;

  //assign uart_0_s1_readyfordata_from_sa = uart_0_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_0_s1_readyfordata_from_sa = uart_0_s1_readyfordata;

  //uart_0_s1_arb_share_counter set values, which is an e_mux
  assign uart_0_s1_arb_share_set_values = (Medipix_sopc_burst_11_downstream_granted_uart_0_s1)? Medipix_sopc_burst_11_downstream_arbitrationshare :
    1;

  //uart_0_s1_non_bursting_master_requests mux, which is an e_mux
  assign uart_0_s1_non_bursting_master_requests = 0;

  //uart_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign uart_0_s1_any_bursting_master_saved_grant = Medipix_sopc_burst_11_downstream_saved_grant_uart_0_s1;

  //uart_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign uart_0_s1_arb_share_counter_next_value = uart_0_s1_firsttransfer ? (uart_0_s1_arb_share_set_values - 1) : |uart_0_s1_arb_share_counter ? (uart_0_s1_arb_share_counter - 1) : 0;

  //uart_0_s1_allgrants all slave grants, which is an e_mux
  assign uart_0_s1_allgrants = |uart_0_s1_grant_vector;

  //uart_0_s1_end_xfer assignment, which is an e_assign
  assign uart_0_s1_end_xfer = ~(uart_0_s1_waits_for_read | uart_0_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_uart_0_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_uart_0_s1 = uart_0_s1_end_xfer & (~uart_0_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //uart_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign uart_0_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_uart_0_s1 & uart_0_s1_allgrants) | (end_xfer_arb_share_counter_term_uart_0_s1 & ~uart_0_s1_non_bursting_master_requests);

  //uart_0_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          uart_0_s1_arb_share_counter <= 0;
      else if (uart_0_s1_arb_counter_enable)
          uart_0_s1_arb_share_counter <= uart_0_s1_arb_share_counter_next_value;
    end


  //uart_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          uart_0_s1_slavearbiterlockenable <= 0;
      else if ((|uart_0_s1_master_qreq_vector & end_xfer_arb_share_counter_term_uart_0_s1) | (end_xfer_arb_share_counter_term_uart_0_s1 & ~uart_0_s1_non_bursting_master_requests))
          uart_0_s1_slavearbiterlockenable <= |uart_0_s1_arb_share_counter_next_value;
    end


  //Medipix_sopc_burst_11/downstream uart_0/s1 arbiterlock, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_arbiterlock = uart_0_s1_slavearbiterlockenable & Medipix_sopc_burst_11_downstream_continuerequest;

  //uart_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign uart_0_s1_slavearbiterlockenable2 = |uart_0_s1_arb_share_counter_next_value;

  //Medipix_sopc_burst_11/downstream uart_0/s1 arbiterlock2, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_arbiterlock2 = uart_0_s1_slavearbiterlockenable2 & Medipix_sopc_burst_11_downstream_continuerequest;

  //uart_0_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign uart_0_s1_any_continuerequest = 1;

  //Medipix_sopc_burst_11_downstream_continuerequest continued request, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_continuerequest = 1;

  assign Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1 = Medipix_sopc_burst_11_downstream_requests_uart_0_s1 & ~((Medipix_sopc_burst_11_downstream_read & ((Medipix_sopc_burst_11_downstream_latency_counter != 0))));
  //local readdatavalid Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1, which is an e_mux
  assign Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1 = Medipix_sopc_burst_11_downstream_granted_uart_0_s1 & Medipix_sopc_burst_11_downstream_read & ~uart_0_s1_waits_for_read;

  //uart_0_s1_writedata mux, which is an e_mux
  assign uart_0_s1_writedata = Medipix_sopc_burst_11_downstream_writedata;

  //master is always granted when requested
  assign Medipix_sopc_burst_11_downstream_granted_uart_0_s1 = Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1;

  //Medipix_sopc_burst_11/downstream saved-grant uart_0/s1, which is an e_assign
  assign Medipix_sopc_burst_11_downstream_saved_grant_uart_0_s1 = Medipix_sopc_burst_11_downstream_requests_uart_0_s1;

  //allow new arb cycle for uart_0/s1, which is an e_assign
  assign uart_0_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign uart_0_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign uart_0_s1_master_qreq_vector = 1;

  assign uart_0_s1_begintransfer = uart_0_s1_begins_xfer;
  //uart_0_s1_reset_n assignment, which is an e_assign
  assign uart_0_s1_reset_n = reset_n;

  assign uart_0_s1_chipselect = Medipix_sopc_burst_11_downstream_granted_uart_0_s1;
  //uart_0_s1_firsttransfer first transaction, which is an e_assign
  assign uart_0_s1_firsttransfer = uart_0_s1_begins_xfer ? uart_0_s1_unreg_firsttransfer : uart_0_s1_reg_firsttransfer;

  //uart_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign uart_0_s1_unreg_firsttransfer = ~(uart_0_s1_slavearbiterlockenable & uart_0_s1_any_continuerequest);

  //uart_0_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          uart_0_s1_reg_firsttransfer <= 1'b1;
      else if (uart_0_s1_begins_xfer)
          uart_0_s1_reg_firsttransfer <= uart_0_s1_unreg_firsttransfer;
    end


  //uart_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign uart_0_s1_beginbursttransfer_internal = uart_0_s1_begins_xfer;

  //~uart_0_s1_read_n assignment, which is an e_mux
  assign uart_0_s1_read_n = ~(Medipix_sopc_burst_11_downstream_granted_uart_0_s1 & Medipix_sopc_burst_11_downstream_read);

  //~uart_0_s1_write_n assignment, which is an e_mux
  assign uart_0_s1_write_n = ~(Medipix_sopc_burst_11_downstream_granted_uart_0_s1 & Medipix_sopc_burst_11_downstream_write);

  //uart_0_s1_address mux, which is an e_mux
  assign uart_0_s1_address = Medipix_sopc_burst_11_downstream_nativeaddress;

  //d1_uart_0_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_uart_0_s1_end_xfer <= 1;
      else 
        d1_uart_0_s1_end_xfer <= uart_0_s1_end_xfer;
    end


  //uart_0_s1_waits_for_read in a cycle, which is an e_mux
  assign uart_0_s1_waits_for_read = uart_0_s1_in_a_read_cycle & uart_0_s1_begins_xfer;

  //uart_0_s1_in_a_read_cycle assignment, which is an e_assign
  assign uart_0_s1_in_a_read_cycle = Medipix_sopc_burst_11_downstream_granted_uart_0_s1 & Medipix_sopc_burst_11_downstream_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = uart_0_s1_in_a_read_cycle;

  //uart_0_s1_waits_for_write in a cycle, which is an e_mux
  assign uart_0_s1_waits_for_write = uart_0_s1_in_a_write_cycle & uart_0_s1_begins_xfer;

  //uart_0_s1_in_a_write_cycle assignment, which is an e_assign
  assign uart_0_s1_in_a_write_cycle = Medipix_sopc_burst_11_downstream_granted_uart_0_s1 & Medipix_sopc_burst_11_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = uart_0_s1_in_a_write_cycle;

  assign wait_for_uart_0_s1_counter = 0;
  //assign uart_0_s1_irq_from_sa = uart_0_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_0_s1_irq_from_sa = uart_0_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //uart_0/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //Medipix_sopc_burst_11/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_11_downstream_requests_uart_0_s1 && (Medipix_sopc_burst_11_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_11/downstream drove 0 on its 'arbitrationshare' port while accessing slave uart_0/s1", $time);
          $stop;
        end
    end


  //Medipix_sopc_burst_11/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (Medipix_sopc_burst_11_downstream_requests_uart_0_s1 && (Medipix_sopc_burst_11_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: Medipix_sopc_burst_11/downstream drove 0 on its 'burstcount' port while accessing slave uart_0/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_reset_ram_aux_half_rate_clk_out_domain_synch_module (
                                                                          // inputs:
                                                                           clk,
                                                                           data_in,
                                                                           reset_n,

                                                                          // outputs:
                                                                           data_out
                                                                        )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc_reset_ram_phy_clk_out_domain_synch_module (
                                                                // inputs:
                                                                 clk,
                                                                 data_in,
                                                                 reset_n,

                                                                // outputs:
                                                                 data_out
                                                              )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Medipix_sopc (
                      // 1) global signals:
                       clk_125,
                       ram_aux_full_rate_clk_out,
                       ram_aux_half_rate_clk_out,
                       ram_phy_clk_out,
                       reset_n,

                      // the_epcs_controller
                       data0_to_the_epcs_controller,
                       dclk_from_the_epcs_controller,
                       sce_from_the_epcs_controller,
                       sdo_from_the_epcs_controller,

                      // the_igor_mac
                       mcoll_pad_i_to_the_igor_mac,
                       mcrs_pad_i_to_the_igor_mac,
                       md_pad_i_to_the_igor_mac,
                       md_pad_o_from_the_igor_mac,
                       md_padoe_o_from_the_igor_mac,
                       mdc_pad_o_from_the_igor_mac,
                       mrx_clk_pad_i_to_the_igor_mac,
                       mrxd_pad_i_to_the_igor_mac,
                       mrxdv_pad_i_to_the_igor_mac,
                       mrxerr_pad_i_to_the_igor_mac,
                       mtx_clk_pad_i_to_the_igor_mac,
                       mtxd_pad_o_from_the_igor_mac,
                       mtxen_pad_o_from_the_igor_mac,
                       mtxerr_pad_o_from_the_igor_mac,

                      // the_ram
                       global_reset_n_to_the_ram,
                       local_init_done_from_the_ram,
                       local_refresh_ack_from_the_ram,
                       local_wdata_req_from_the_ram,
                       mem_addr_from_the_ram,
                       mem_ba_from_the_ram,
                       mem_cas_n_from_the_ram,
                       mem_cke_from_the_ram,
                       mem_clk_n_to_and_from_the_ram,
                       mem_clk_to_and_from_the_ram,
                       mem_cs_n_from_the_ram,
                       mem_dm_from_the_ram,
                       mem_dq_to_and_from_the_ram,
                       mem_dqs_to_and_from_the_ram,
                       mem_odt_from_the_ram,
                       mem_ras_n_from_the_ram,
                       mem_we_n_from_the_ram,
                       reset_phy_clk_n_from_the_ram,

                      // the_spi_0
                       MISO_to_the_spi_0,
                       MOSI_from_the_spi_0,
                       SCLK_from_the_spi_0,
                       SS_n_from_the_spi_0,

                      // the_tx_table
                       clock_vhdl_to_the_tx_table,
                       in_Nreset_to_the_tx_table,
                       info_out_from_the_tx_table,
                       irq_from_the_tx_table,
                       out_data_from_the_tx_table,
                       out_sync_from_the_tx_table,
                       out_valid_from_the_tx_table,

                      // the_uart_0
                       rxd_to_the_uart_0,
                       txd_from_the_uart_0
                    )
;

  output           MOSI_from_the_spi_0;
  output           SCLK_from_the_spi_0;
  output  [  1: 0] SS_n_from_the_spi_0;
  output           dclk_from_the_epcs_controller;
  output  [  7: 0] info_out_from_the_tx_table;
  output           irq_from_the_tx_table;
  output           local_init_done_from_the_ram;
  output           local_refresh_ack_from_the_ram;
  output           local_wdata_req_from_the_ram;
  output           md_pad_o_from_the_igor_mac;
  output           md_padoe_o_from_the_igor_mac;
  output           mdc_pad_o_from_the_igor_mac;
  output  [ 12: 0] mem_addr_from_the_ram;
  output  [  2: 0] mem_ba_from_the_ram;
  output           mem_cas_n_from_the_ram;
  output           mem_cke_from_the_ram;
  inout            mem_clk_n_to_and_from_the_ram;
  inout            mem_clk_to_and_from_the_ram;
  output           mem_cs_n_from_the_ram;
  output  [  1: 0] mem_dm_from_the_ram;
  inout   [ 15: 0] mem_dq_to_and_from_the_ram;
  inout   [  1: 0] mem_dqs_to_and_from_the_ram;
  output           mem_odt_from_the_ram;
  output           mem_ras_n_from_the_ram;
  output           mem_we_n_from_the_ram;
  output  [  3: 0] mtxd_pad_o_from_the_igor_mac;
  output           mtxen_pad_o_from_the_igor_mac;
  output           mtxerr_pad_o_from_the_igor_mac;
  output  [  7: 0] out_data_from_the_tx_table;
  output           out_sync_from_the_tx_table;
  output           out_valid_from_the_tx_table;
  output           ram_aux_full_rate_clk_out;
  output           ram_aux_half_rate_clk_out;
  output           ram_phy_clk_out;
  output           reset_phy_clk_n_from_the_ram;
  output           sce_from_the_epcs_controller;
  output           sdo_from_the_epcs_controller;
  output           txd_from_the_uart_0;
  input            MISO_to_the_spi_0;
  input            clk_125;
  input            clock_vhdl_to_the_tx_table;
  input            data0_to_the_epcs_controller;
  input            global_reset_n_to_the_ram;
  input            in_Nreset_to_the_tx_table;
  input            mcoll_pad_i_to_the_igor_mac;
  input            mcrs_pad_i_to_the_igor_mac;
  input            md_pad_i_to_the_igor_mac;
  input            mrx_clk_pad_i_to_the_igor_mac;
  input   [  3: 0] mrxd_pad_i_to_the_igor_mac;
  input            mrxdv_pad_i_to_the_igor_mac;
  input            mrxerr_pad_i_to_the_igor_mac;
  input            mtx_clk_pad_i_to_the_igor_mac;
  input            reset_n;
  input            rxd_to_the_uart_0;

  wire             MOSI_from_the_spi_0;
  wire    [ 10: 0] Medipix_sopc_burst_0_downstream_address;
  wire    [ 10: 0] Medipix_sopc_burst_0_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_0_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_0_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_0_downstream_byteenable;
  wire             Medipix_sopc_burst_0_downstream_debugaccess;
  wire             Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_latency_counter;
  wire    [ 10: 0] Medipix_sopc_burst_0_downstream_nativeaddress;
  wire             Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_read;
  wire             Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  wire    [ 31: 0] Medipix_sopc_burst_0_downstream_readdata;
  wire             Medipix_sopc_burst_0_downstream_readdatavalid;
  wire             Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_0_downstream_reset_n;
  wire             Medipix_sopc_burst_0_downstream_waitrequest;
  wire             Medipix_sopc_burst_0_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_0_downstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_0_upstream_address;
  wire    [ 12: 0] Medipix_sopc_burst_0_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_0_upstream_byteenable;
  wire             Medipix_sopc_burst_0_upstream_debugaccess;
  wire             Medipix_sopc_burst_0_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_0_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_0_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_0_upstream_readdatavalid;
  wire             Medipix_sopc_burst_0_upstream_waitrequest;
  wire             Medipix_sopc_burst_0_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_0_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_0_upstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_10_downstream_address;
  wire    [  3: 0] Medipix_sopc_burst_10_downstream_address_to_slave;
  wire    [  4: 0] Medipix_sopc_burst_10_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_10_downstream_burstcount;
  wire    [  1: 0] Medipix_sopc_burst_10_downstream_byteenable;
  wire             Medipix_sopc_burst_10_downstream_debugaccess;
  wire             Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_latency_counter;
  wire    [  3: 0] Medipix_sopc_burst_10_downstream_nativeaddress;
  wire             Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_read;
  wire             Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port;
  wire    [ 15: 0] Medipix_sopc_burst_10_downstream_readdata;
  wire             Medipix_sopc_burst_10_downstream_readdatavalid;
  wire             Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port;
  wire             Medipix_sopc_burst_10_downstream_reset_n;
  wire             Medipix_sopc_burst_10_downstream_waitrequest;
  wire             Medipix_sopc_burst_10_downstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_10_downstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_10_upstream_burstcount;
  wire    [  4: 0] Medipix_sopc_burst_10_upstream_byteaddress;
  wire    [  1: 0] Medipix_sopc_burst_10_upstream_byteenable;
  wire             Medipix_sopc_burst_10_upstream_debugaccess;
  wire             Medipix_sopc_burst_10_upstream_read;
  wire    [ 15: 0] Medipix_sopc_burst_10_upstream_readdata;
  wire    [ 15: 0] Medipix_sopc_burst_10_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_10_upstream_readdatavalid;
  wire             Medipix_sopc_burst_10_upstream_waitrequest;
  wire             Medipix_sopc_burst_10_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_10_upstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_10_upstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_11_downstream_address;
  wire    [  3: 0] Medipix_sopc_burst_11_downstream_address_to_slave;
  wire    [  4: 0] Medipix_sopc_burst_11_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_11_downstream_burstcount;
  wire    [  1: 0] Medipix_sopc_burst_11_downstream_byteenable;
  wire             Medipix_sopc_burst_11_downstream_debugaccess;
  wire             Medipix_sopc_burst_11_downstream_granted_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_latency_counter;
  wire    [  3: 0] Medipix_sopc_burst_11_downstream_nativeaddress;
  wire             Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_read;
  wire             Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1;
  wire    [ 15: 0] Medipix_sopc_burst_11_downstream_readdata;
  wire             Medipix_sopc_burst_11_downstream_readdatavalid;
  wire             Medipix_sopc_burst_11_downstream_requests_uart_0_s1;
  wire             Medipix_sopc_burst_11_downstream_reset_n;
  wire             Medipix_sopc_burst_11_downstream_waitrequest;
  wire             Medipix_sopc_burst_11_downstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_11_downstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_11_upstream_burstcount;
  wire    [  4: 0] Medipix_sopc_burst_11_upstream_byteaddress;
  wire    [  1: 0] Medipix_sopc_burst_11_upstream_byteenable;
  wire             Medipix_sopc_burst_11_upstream_debugaccess;
  wire             Medipix_sopc_burst_11_upstream_read;
  wire    [ 15: 0] Medipix_sopc_burst_11_upstream_readdata;
  wire    [ 15: 0] Medipix_sopc_burst_11_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_11_upstream_readdatavalid;
  wire             Medipix_sopc_burst_11_upstream_waitrequest;
  wire             Medipix_sopc_burst_11_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_11_upstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_11_upstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_1_downstream_address;
  wire    [ 10: 0] Medipix_sopc_burst_1_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_1_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_1_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_1_downstream_byteenable;
  wire             Medipix_sopc_burst_1_downstream_debugaccess;
  wire             Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_latency_counter;
  wire    [ 10: 0] Medipix_sopc_burst_1_downstream_nativeaddress;
  wire             Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_read;
  wire             Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module;
  wire    [ 31: 0] Medipix_sopc_burst_1_downstream_readdata;
  wire             Medipix_sopc_burst_1_downstream_readdatavalid;
  wire             Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module;
  wire             Medipix_sopc_burst_1_downstream_reset_n;
  wire             Medipix_sopc_burst_1_downstream_waitrequest;
  wire             Medipix_sopc_burst_1_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_1_downstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_1_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_burstcount;
  wire    [ 12: 0] Medipix_sopc_burst_1_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_1_upstream_byteenable;
  wire             Medipix_sopc_burst_1_upstream_debugaccess;
  wire             Medipix_sopc_burst_1_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_1_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_1_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_1_upstream_readdatavalid;
  wire             Medipix_sopc_burst_1_upstream_waitrequest;
  wire             Medipix_sopc_burst_1_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_1_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_1_upstream_writedata;
  wire    [  2: 0] Medipix_sopc_burst_2_downstream_address;
  wire    [  2: 0] Medipix_sopc_burst_2_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_2_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_2_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_2_downstream_byteenable;
  wire             Medipix_sopc_burst_2_downstream_debugaccess;
  wire             Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_latency_counter;
  wire    [  2: 0] Medipix_sopc_burst_2_downstream_nativeaddress;
  wire             Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_read;
  wire             Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  wire    [ 31: 0] Medipix_sopc_burst_2_downstream_readdata;
  wire             Medipix_sopc_burst_2_downstream_readdatavalid;
  wire             Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave;
  wire             Medipix_sopc_burst_2_downstream_reset_n;
  wire             Medipix_sopc_burst_2_downstream_waitrequest;
  wire             Medipix_sopc_burst_2_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_2_downstream_writedata;
  wire    [  2: 0] Medipix_sopc_burst_2_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_burstcount;
  wire    [  4: 0] Medipix_sopc_burst_2_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_2_upstream_byteenable;
  wire             Medipix_sopc_burst_2_upstream_debugaccess;
  wire             Medipix_sopc_burst_2_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_2_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_2_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_2_upstream_readdatavalid;
  wire             Medipix_sopc_burst_2_upstream_waitrequest;
  wire             Medipix_sopc_burst_2_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_2_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_2_upstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_3_downstream_address;
  wire    [  3: 0] Medipix_sopc_burst_3_downstream_address_to_slave;
  wire    [  4: 0] Medipix_sopc_burst_3_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_3_downstream_burstcount;
  wire    [  1: 0] Medipix_sopc_burst_3_downstream_byteenable;
  wire             Medipix_sopc_burst_3_downstream_debugaccess;
  wire             Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_latency_counter;
  wire    [  3: 0] Medipix_sopc_burst_3_downstream_nativeaddress;
  wire             Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_read;
  wire             Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1;
  wire    [ 15: 0] Medipix_sopc_burst_3_downstream_readdata;
  wire             Medipix_sopc_burst_3_downstream_readdatavalid;
  wire             Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1;
  wire             Medipix_sopc_burst_3_downstream_reset_n;
  wire             Medipix_sopc_burst_3_downstream_waitrequest;
  wire             Medipix_sopc_burst_3_downstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_3_downstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_3_upstream_burstcount;
  wire    [  4: 0] Medipix_sopc_burst_3_upstream_byteaddress;
  wire    [  1: 0] Medipix_sopc_burst_3_upstream_byteenable;
  wire             Medipix_sopc_burst_3_upstream_debugaccess;
  wire             Medipix_sopc_burst_3_upstream_read;
  wire    [ 15: 0] Medipix_sopc_burst_3_upstream_readdata;
  wire    [ 15: 0] Medipix_sopc_burst_3_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_3_upstream_readdatavalid;
  wire             Medipix_sopc_burst_3_upstream_waitrequest;
  wire             Medipix_sopc_burst_3_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_3_upstream_write;
  wire    [ 15: 0] Medipix_sopc_burst_3_upstream_writedata;
  wire    [ 26: 0] Medipix_sopc_burst_4_downstream_address;
  wire    [ 26: 0] Medipix_sopc_burst_4_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_4_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_4_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_4_downstream_byteenable;
  wire             Medipix_sopc_burst_4_downstream_debugaccess;
  wire             Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_latency_counter;
  wire    [ 26: 0] Medipix_sopc_burst_4_downstream_nativeaddress;
  wire             Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_read;
  wire             Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register;
  wire    [ 31: 0] Medipix_sopc_burst_4_downstream_readdata;
  wire             Medipix_sopc_burst_4_downstream_readdatavalid;
  wire             Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1;
  wire             Medipix_sopc_burst_4_downstream_reset_n;
  wire             Medipix_sopc_burst_4_downstream_waitrequest;
  wire             Medipix_sopc_burst_4_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_4_downstream_writedata;
  wire    [ 26: 0] Medipix_sopc_burst_4_upstream_address;
  wire    [ 28: 0] Medipix_sopc_burst_4_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_4_upstream_byteenable;
  wire             Medipix_sopc_burst_4_upstream_debugaccess;
  wire             Medipix_sopc_burst_4_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_4_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_4_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_4_upstream_readdatavalid;
  wire             Medipix_sopc_burst_4_upstream_waitrequest;
  wire             Medipix_sopc_burst_4_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_4_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_4_upstream_writedata;
  wire    [ 26: 0] Medipix_sopc_burst_5_downstream_address;
  wire    [ 26: 0] Medipix_sopc_burst_5_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_5_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_5_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_5_downstream_byteenable;
  wire             Medipix_sopc_burst_5_downstream_debugaccess;
  wire             Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_latency_counter;
  wire    [ 26: 0] Medipix_sopc_burst_5_downstream_nativeaddress;
  wire             Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_read;
  wire             Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register;
  wire    [ 31: 0] Medipix_sopc_burst_5_downstream_readdata;
  wire             Medipix_sopc_burst_5_downstream_readdatavalid;
  wire             Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1;
  wire             Medipix_sopc_burst_5_downstream_reset_n;
  wire             Medipix_sopc_burst_5_downstream_waitrequest;
  wire             Medipix_sopc_burst_5_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_5_downstream_writedata;
  wire    [ 26: 0] Medipix_sopc_burst_5_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_burstcount;
  wire    [ 28: 0] Medipix_sopc_burst_5_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_5_upstream_byteenable;
  wire             Medipix_sopc_burst_5_upstream_debugaccess;
  wire             Medipix_sopc_burst_5_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_5_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_5_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_5_upstream_readdatavalid;
  wire             Medipix_sopc_burst_5_upstream_waitrequest;
  wire             Medipix_sopc_burst_5_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_5_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_5_upstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_6_downstream_address;
  wire    [ 10: 0] Medipix_sopc_burst_6_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_6_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_6_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_6_downstream_byteenable;
  wire             Medipix_sopc_burst_6_downstream_debugaccess;
  wire             Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_latency_counter;
  wire    [ 10: 0] Medipix_sopc_burst_6_downstream_nativeaddress;
  wire             Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_read;
  wire             Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port;
  wire    [ 31: 0] Medipix_sopc_burst_6_downstream_readdata;
  wire             Medipix_sopc_burst_6_downstream_readdatavalid;
  wire             Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_6_downstream_reset_n;
  wire             Medipix_sopc_burst_6_downstream_waitrequest;
  wire             Medipix_sopc_burst_6_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_6_downstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_6_upstream_address;
  wire    [ 12: 0] Medipix_sopc_burst_6_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_6_upstream_byteenable;
  wire             Medipix_sopc_burst_6_upstream_debugaccess;
  wire             Medipix_sopc_burst_6_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_6_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_6_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_6_upstream_readdatavalid;
  wire             Medipix_sopc_burst_6_upstream_waitrequest;
  wire             Medipix_sopc_burst_6_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_6_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_6_upstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_7_downstream_address;
  wire    [ 10: 0] Medipix_sopc_burst_7_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_7_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_7_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_7_downstream_byteenable;
  wire             Medipix_sopc_burst_7_downstream_debugaccess;
  wire             Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_latency_counter;
  wire    [ 10: 0] Medipix_sopc_burst_7_downstream_nativeaddress;
  wire             Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_read;
  wire             Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port;
  wire    [ 31: 0] Medipix_sopc_burst_7_downstream_readdata;
  wire             Medipix_sopc_burst_7_downstream_readdatavalid;
  wire             Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port;
  wire             Medipix_sopc_burst_7_downstream_reset_n;
  wire             Medipix_sopc_burst_7_downstream_waitrequest;
  wire             Medipix_sopc_burst_7_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_7_downstream_writedata;
  wire    [ 10: 0] Medipix_sopc_burst_7_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_burstcount;
  wire    [ 12: 0] Medipix_sopc_burst_7_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_7_upstream_byteenable;
  wire             Medipix_sopc_burst_7_upstream_debugaccess;
  wire             Medipix_sopc_burst_7_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_7_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_7_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_7_upstream_readdatavalid;
  wire             Medipix_sopc_burst_7_upstream_waitrequest;
  wire             Medipix_sopc_burst_7_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_7_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_7_upstream_writedata;
  wire    [ 11: 0] Medipix_sopc_burst_8_downstream_address;
  wire    [ 11: 0] Medipix_sopc_burst_8_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_8_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_8_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_8_downstream_byteenable;
  wire             Medipix_sopc_burst_8_downstream_debugaccess;
  wire             Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_latency_counter;
  wire    [ 11: 0] Medipix_sopc_burst_8_downstream_nativeaddress;
  wire             Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_read;
  wire             Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port;
  wire    [ 31: 0] Medipix_sopc_burst_8_downstream_readdata;
  wire             Medipix_sopc_burst_8_downstream_readdatavalid;
  wire             Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port;
  wire             Medipix_sopc_burst_8_downstream_reset_n;
  wire             Medipix_sopc_burst_8_downstream_waitrequest;
  wire             Medipix_sopc_burst_8_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_8_downstream_writedata;
  wire    [ 11: 0] Medipix_sopc_burst_8_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_burstcount;
  wire    [ 13: 0] Medipix_sopc_burst_8_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_8_upstream_byteenable;
  wire             Medipix_sopc_burst_8_upstream_debugaccess;
  wire             Medipix_sopc_burst_8_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_8_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_8_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_8_upstream_readdatavalid;
  wire             Medipix_sopc_burst_8_upstream_waitrequest;
  wire             Medipix_sopc_burst_8_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_8_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_8_upstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_address;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_address_to_slave;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_arbitrationshare;
  wire             Medipix_sopc_burst_9_downstream_burstcount;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_byteenable;
  wire             Medipix_sopc_burst_9_downstream_debugaccess;
  wire             Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_latency_counter;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_nativeaddress;
  wire             Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_read;
  wire             Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0;
  wire    [ 31: 0] Medipix_sopc_burst_9_downstream_readdata;
  wire             Medipix_sopc_burst_9_downstream_readdatavalid;
  wire             Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0;
  wire             Medipix_sopc_burst_9_downstream_reset_n;
  wire             Medipix_sopc_burst_9_downstream_waitrequest;
  wire             Medipix_sopc_burst_9_downstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_9_downstream_writedata;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_address;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_burstcount;
  wire    [  5: 0] Medipix_sopc_burst_9_upstream_byteaddress;
  wire    [  3: 0] Medipix_sopc_burst_9_upstream_byteenable;
  wire             Medipix_sopc_burst_9_upstream_debugaccess;
  wire             Medipix_sopc_burst_9_upstream_read;
  wire    [ 31: 0] Medipix_sopc_burst_9_upstream_readdata;
  wire    [ 31: 0] Medipix_sopc_burst_9_upstream_readdata_from_sa;
  wire             Medipix_sopc_burst_9_upstream_readdatavalid;
  wire             Medipix_sopc_burst_9_upstream_waitrequest;
  wire             Medipix_sopc_burst_9_upstream_waitrequest_from_sa;
  wire             Medipix_sopc_burst_9_upstream_write;
  wire    [ 31: 0] Medipix_sopc_burst_9_upstream_writedata;
  wire             SCLK_from_the_spi_0;
  wire    [  1: 0] SS_n_from_the_spi_0;
  wire             clk_125_reset_n;
  wire    [ 26: 0] clock_crossing_m1_address;
  wire    [ 26: 0] clock_crossing_m1_address_to_slave;
  wire    [  3: 0] clock_crossing_m1_byteenable;
  wire             clock_crossing_m1_endofpacket;
  wire             clock_crossing_m1_granted_ram_s1;
  wire             clock_crossing_m1_latency_counter;
  wire    [ 24: 0] clock_crossing_m1_nativeaddress;
  wire             clock_crossing_m1_qualified_request_ram_s1;
  wire             clock_crossing_m1_read;
  wire             clock_crossing_m1_read_data_valid_ram_s1;
  wire             clock_crossing_m1_read_data_valid_ram_s1_shift_register;
  wire    [ 31: 0] clock_crossing_m1_readdata;
  wire             clock_crossing_m1_readdatavalid;
  wire             clock_crossing_m1_requests_ram_s1;
  wire             clock_crossing_m1_reset_n;
  wire             clock_crossing_m1_waitrequest;
  wire             clock_crossing_m1_write;
  wire    [ 31: 0] clock_crossing_m1_writedata;
  wire    [ 24: 0] clock_crossing_s1_address;
  wire    [  3: 0] clock_crossing_s1_byteenable;
  wire             clock_crossing_s1_endofpacket;
  wire             clock_crossing_s1_endofpacket_from_sa;
  wire    [ 24: 0] clock_crossing_s1_nativeaddress;
  wire             clock_crossing_s1_read;
  wire    [ 31: 0] clock_crossing_s1_readdata;
  wire    [ 31: 0] clock_crossing_s1_readdata_from_sa;
  wire             clock_crossing_s1_readdatavalid;
  wire             clock_crossing_s1_reset_n;
  wire             clock_crossing_s1_waitrequest;
  wire             clock_crossing_s1_waitrequest_from_sa;
  wire             clock_crossing_s1_write;
  wire    [ 31: 0] clock_crossing_s1_writedata;
  wire    [ 27: 0] cpu_linux_data_master_address;
  wire    [ 27: 0] cpu_linux_data_master_address_to_slave;
  wire    [  3: 0] cpu_linux_data_master_burstcount;
  wire    [  3: 0] cpu_linux_data_master_byteenable;
  wire             cpu_linux_data_master_debugaccess;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream;
  wire    [ 31: 0] cpu_linux_data_master_irq;
  wire             cpu_linux_data_master_latency_counter;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_read;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register;
  wire    [ 31: 0] cpu_linux_data_master_readdata;
  wire             cpu_linux_data_master_readdatavalid;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream;
  wire             cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream;
  wire             cpu_linux_data_master_waitrequest;
  wire             cpu_linux_data_master_write;
  wire    [ 31: 0] cpu_linux_data_master_writedata;
  wire    [ 27: 0] cpu_linux_instruction_master_address;
  wire    [ 27: 0] cpu_linux_instruction_master_address_to_slave;
  wire    [  3: 0] cpu_linux_instruction_master_burstcount;
  wire             cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_latency_counter;
  wire             cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_read;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register;
  wire    [ 31: 0] cpu_linux_instruction_master_readdata;
  wire             cpu_linux_instruction_master_readdatavalid;
  wire             cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream;
  wire             cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream;
  wire             cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream;
  wire             cpu_linux_instruction_master_waitrequest;
  wire    [  8: 0] cpu_linux_jtag_debug_module_address;
  wire             cpu_linux_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_linux_jtag_debug_module_byteenable;
  wire             cpu_linux_jtag_debug_module_chipselect;
  wire             cpu_linux_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_linux_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_linux_jtag_debug_module_readdata_from_sa;
  wire             cpu_linux_jtag_debug_module_reset_n;
  wire             cpu_linux_jtag_debug_module_resetrequest;
  wire             cpu_linux_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_linux_jtag_debug_module_write;
  wire    [ 31: 0] cpu_linux_jtag_debug_module_writedata;
  wire             d1_Medipix_sopc_burst_0_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_10_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_11_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_1_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_2_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_3_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_4_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_5_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_6_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_7_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_8_upstream_end_xfer;
  wire             d1_Medipix_sopc_burst_9_upstream_end_xfer;
  wire             d1_clock_crossing_s1_end_xfer;
  wire             d1_cpu_linux_jtag_debug_module_end_xfer;
  wire             d1_epcs_controller_epcs_control_port_end_xfer;
  wire             d1_igor_mac_control_port_end_xfer;
  wire             d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  wire             d1_ram_s1_end_xfer;
  wire             d1_spi_0_spi_control_port_end_xfer;
  wire             d1_sys_clk_freq_s1_end_xfer;
  wire             d1_tx_table_avalon_slave_0_end_xfer;
  wire             d1_uart_0_s1_end_xfer;
  wire             dclk_from_the_epcs_controller;
  wire    [  8: 0] epcs_controller_epcs_control_port_address;
  wire             epcs_controller_epcs_control_port_chipselect;
  wire             epcs_controller_epcs_control_port_dataavailable;
  wire             epcs_controller_epcs_control_port_dataavailable_from_sa;
  wire             epcs_controller_epcs_control_port_endofpacket;
  wire             epcs_controller_epcs_control_port_endofpacket_from_sa;
  wire             epcs_controller_epcs_control_port_irq;
  wire             epcs_controller_epcs_control_port_irq_from_sa;
  wire             epcs_controller_epcs_control_port_read_n;
  wire    [ 31: 0] epcs_controller_epcs_control_port_readdata;
  wire    [ 31: 0] epcs_controller_epcs_control_port_readdata_from_sa;
  wire             epcs_controller_epcs_control_port_readyfordata;
  wire             epcs_controller_epcs_control_port_readyfordata_from_sa;
  wire             epcs_controller_epcs_control_port_reset_n;
  wire             epcs_controller_epcs_control_port_write_n;
  wire    [ 31: 0] epcs_controller_epcs_control_port_writedata;
  wire    [  9: 0] igor_mac_control_port_address;
  wire             igor_mac_control_port_chipselect;
  wire             igor_mac_control_port_irq;
  wire             igor_mac_control_port_irq_from_sa;
  wire             igor_mac_control_port_read;
  wire    [ 31: 0] igor_mac_control_port_readdata;
  wire    [ 31: 0] igor_mac_control_port_readdata_from_sa;
  wire             igor_mac_control_port_reset;
  wire             igor_mac_control_port_waitrequest_n;
  wire             igor_mac_control_port_waitrequest_n_from_sa;
  wire             igor_mac_control_port_write;
  wire    [ 31: 0] igor_mac_control_port_writedata;
  wire    [ 31: 0] igor_mac_rx_master_address;
  wire    [ 31: 0] igor_mac_rx_master_address_to_slave;
  wire    [  3: 0] igor_mac_rx_master_byteenable;
  wire             igor_mac_rx_master_granted_clock_crossing_s1;
  wire             igor_mac_rx_master_qualified_request_clock_crossing_s1;
  wire             igor_mac_rx_master_requests_clock_crossing_s1;
  wire             igor_mac_rx_master_waitrequest;
  wire             igor_mac_rx_master_write;
  wire    [ 31: 0] igor_mac_rx_master_writedata;
  wire    [ 31: 0] igor_mac_tx_master_address;
  wire    [ 31: 0] igor_mac_tx_master_address_to_slave;
  wire             igor_mac_tx_master_granted_clock_crossing_s1;
  wire             igor_mac_tx_master_latency_counter;
  wire             igor_mac_tx_master_qualified_request_clock_crossing_s1;
  wire             igor_mac_tx_master_read;
  wire             igor_mac_tx_master_read_data_valid_clock_crossing_s1;
  wire             igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register;
  wire    [ 31: 0] igor_mac_tx_master_readdata;
  wire             igor_mac_tx_master_readdatavalid;
  wire             igor_mac_tx_master_requests_clock_crossing_s1;
  wire             igor_mac_tx_master_waitrequest;
  wire    [  7: 0] info_out_from_the_tx_table;
  wire             irq_from_the_tx_table;
  wire             jtag_uart_0_avalon_jtag_slave_address;
  wire             jtag_uart_0_avalon_jtag_slave_chipselect;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_irq;
  wire             jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_reset_n;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  wire             local_init_done_from_the_ram;
  wire             local_refresh_ack_from_the_ram;
  wire             local_wdata_req_from_the_ram;
  wire             md_pad_o_from_the_igor_mac;
  wire             md_padoe_o_from_the_igor_mac;
  wire             mdc_pad_o_from_the_igor_mac;
  wire    [ 12: 0] mem_addr_from_the_ram;
  wire    [  2: 0] mem_ba_from_the_ram;
  wire             mem_cas_n_from_the_ram;
  wire             mem_cke_from_the_ram;
  wire             mem_clk_n_to_and_from_the_ram;
  wire             mem_clk_to_and_from_the_ram;
  wire             mem_cs_n_from_the_ram;
  wire    [  1: 0] mem_dm_from_the_ram;
  wire    [ 15: 0] mem_dq_to_and_from_the_ram;
  wire    [  1: 0] mem_dqs_to_and_from_the_ram;
  wire             mem_odt_from_the_ram;
  wire             mem_ras_n_from_the_ram;
  wire             mem_we_n_from_the_ram;
  wire    [  3: 0] mtxd_pad_o_from_the_igor_mac;
  wire             mtxen_pad_o_from_the_igor_mac;
  wire             mtxerr_pad_o_from_the_igor_mac;
  wire             out_clk_ram_aux_full_rate_clk;
  wire             out_clk_ram_aux_half_rate_clk;
  wire             out_clk_ram_phy_clk;
  wire    [  7: 0] out_data_from_the_tx_table;
  wire             out_sync_from_the_tx_table;
  wire             out_valid_from_the_tx_table;
  wire             ram_aux_full_rate_clk_out;
  wire             ram_aux_half_rate_clk_out;
  wire             ram_aux_half_rate_clk_out_reset_n;
  wire             ram_phy_clk_out;
  wire             ram_phy_clk_out_reset_n;
  wire    [ 24: 0] ram_s1_address;
  wire             ram_s1_beginbursttransfer;
  wire    [  2: 0] ram_s1_burstcount;
  wire    [  3: 0] ram_s1_byteenable;
  wire             ram_s1_read;
  wire    [ 31: 0] ram_s1_readdata;
  wire    [ 31: 0] ram_s1_readdata_from_sa;
  wire             ram_s1_readdatavalid;
  wire             ram_s1_resetrequest_n;
  wire             ram_s1_resetrequest_n_from_sa;
  wire             ram_s1_waitrequest_n;
  wire             ram_s1_waitrequest_n_from_sa;
  wire             ram_s1_write;
  wire    [ 31: 0] ram_s1_writedata;
  wire             reset_n_sources;
  wire             reset_phy_clk_n_from_the_ram;
  wire             sce_from_the_epcs_controller;
  wire             sdo_from_the_epcs_controller;
  wire    [  2: 0] spi_0_spi_control_port_address;
  wire             spi_0_spi_control_port_chipselect;
  wire             spi_0_spi_control_port_dataavailable;
  wire             spi_0_spi_control_port_dataavailable_from_sa;
  wire             spi_0_spi_control_port_endofpacket;
  wire             spi_0_spi_control_port_endofpacket_from_sa;
  wire             spi_0_spi_control_port_irq;
  wire             spi_0_spi_control_port_irq_from_sa;
  wire             spi_0_spi_control_port_read_n;
  wire    [ 15: 0] spi_0_spi_control_port_readdata;
  wire    [ 15: 0] spi_0_spi_control_port_readdata_from_sa;
  wire             spi_0_spi_control_port_readyfordata;
  wire             spi_0_spi_control_port_readyfordata_from_sa;
  wire             spi_0_spi_control_port_reset_n;
  wire             spi_0_spi_control_port_write_n;
  wire    [ 15: 0] spi_0_spi_control_port_writedata;
  wire    [  2: 0] sys_clk_freq_s1_address;
  wire             sys_clk_freq_s1_chipselect;
  wire             sys_clk_freq_s1_irq;
  wire             sys_clk_freq_s1_irq_from_sa;
  wire    [ 15: 0] sys_clk_freq_s1_readdata;
  wire    [ 15: 0] sys_clk_freq_s1_readdata_from_sa;
  wire             sys_clk_freq_s1_reset_n;
  wire             sys_clk_freq_s1_write_n;
  wire    [ 15: 0] sys_clk_freq_s1_writedata;
  wire    [  1: 0] tx_table_avalon_slave_0_address;
  wire             tx_table_avalon_slave_0_chipselect;
  wire             tx_table_avalon_slave_0_read;
  wire    [ 31: 0] tx_table_avalon_slave_0_readdata;
  wire    [ 31: 0] tx_table_avalon_slave_0_readdata_from_sa;
  wire             tx_table_avalon_slave_0_reset_n;
  wire             tx_table_avalon_slave_0_write;
  wire    [ 31: 0] tx_table_avalon_slave_0_writedata;
  wire             txd_from_the_uart_0;
  wire    [  2: 0] uart_0_s1_address;
  wire             uart_0_s1_begintransfer;
  wire             uart_0_s1_chipselect;
  wire             uart_0_s1_dataavailable;
  wire             uart_0_s1_dataavailable_from_sa;
  wire             uart_0_s1_irq;
  wire             uart_0_s1_irq_from_sa;
  wire             uart_0_s1_read_n;
  wire    [ 15: 0] uart_0_s1_readdata;
  wire    [ 15: 0] uart_0_s1_readdata_from_sa;
  wire             uart_0_s1_readyfordata;
  wire             uart_0_s1_readyfordata_from_sa;
  wire             uart_0_s1_reset_n;
  wire             uart_0_s1_write_n;
  wire    [ 15: 0] uart_0_s1_writedata;
  Medipix_sopc_burst_0_upstream_arbitrator the_Medipix_sopc_burst_0_upstream
    (
      .Medipix_sopc_burst_0_upstream_address                                                     (Medipix_sopc_burst_0_upstream_address),
      .Medipix_sopc_burst_0_upstream_byteaddress                                                 (Medipix_sopc_burst_0_upstream_byteaddress),
      .Medipix_sopc_burst_0_upstream_byteenable                                                  (Medipix_sopc_burst_0_upstream_byteenable),
      .Medipix_sopc_burst_0_upstream_debugaccess                                                 (Medipix_sopc_burst_0_upstream_debugaccess),
      .Medipix_sopc_burst_0_upstream_read                                                        (Medipix_sopc_burst_0_upstream_read),
      .Medipix_sopc_burst_0_upstream_readdata                                                    (Medipix_sopc_burst_0_upstream_readdata),
      .Medipix_sopc_burst_0_upstream_readdata_from_sa                                            (Medipix_sopc_burst_0_upstream_readdata_from_sa),
      .Medipix_sopc_burst_0_upstream_readdatavalid                                               (Medipix_sopc_burst_0_upstream_readdatavalid),
      .Medipix_sopc_burst_0_upstream_waitrequest                                                 (Medipix_sopc_burst_0_upstream_waitrequest),
      .Medipix_sopc_burst_0_upstream_waitrequest_from_sa                                         (Medipix_sopc_burst_0_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_0_upstream_write                                                       (Medipix_sopc_burst_0_upstream_write),
      .clk                                                                                       (ram_aux_half_rate_clk_out),
      .cpu_linux_instruction_master_address_to_slave                                             (cpu_linux_instruction_master_address_to_slave),
      .cpu_linux_instruction_master_burstcount                                                   (cpu_linux_instruction_master_burstcount),
      .cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream                        (cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_latency_counter                                              (cpu_linux_instruction_master_latency_counter),
      .cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream              (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_read                                                         (cpu_linux_instruction_master_read),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream                (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register),
      .cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream                       (cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream),
      .d1_Medipix_sopc_burst_0_upstream_end_xfer                                                 (d1_Medipix_sopc_burst_0_upstream_end_xfer),
      .reset_n                                                                                   (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_0_downstream_arbitrator the_Medipix_sopc_burst_0_downstream
    (
      .Medipix_sopc_burst_0_downstream_address                                       (Medipix_sopc_burst_0_downstream_address),
      .Medipix_sopc_burst_0_downstream_address_to_slave                              (Medipix_sopc_burst_0_downstream_address_to_slave),
      .Medipix_sopc_burst_0_downstream_burstcount                                    (Medipix_sopc_burst_0_downstream_burstcount),
      .Medipix_sopc_burst_0_downstream_byteenable                                    (Medipix_sopc_burst_0_downstream_byteenable),
      .Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module           (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_latency_counter                               (Medipix_sopc_burst_0_downstream_latency_counter),
      .Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module (Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_read                                          (Medipix_sopc_burst_0_downstream_read),
      .Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module   (Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_readdata                                      (Medipix_sopc_burst_0_downstream_readdata),
      .Medipix_sopc_burst_0_downstream_readdatavalid                                 (Medipix_sopc_burst_0_downstream_readdatavalid),
      .Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module          (Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_reset_n                                       (Medipix_sopc_burst_0_downstream_reset_n),
      .Medipix_sopc_burst_0_downstream_waitrequest                                   (Medipix_sopc_burst_0_downstream_waitrequest),
      .Medipix_sopc_burst_0_downstream_write                                         (Medipix_sopc_burst_0_downstream_write),
      .Medipix_sopc_burst_0_downstream_writedata                                     (Medipix_sopc_burst_0_downstream_writedata),
      .clk                                                                           (ram_aux_half_rate_clk_out),
      .cpu_linux_jtag_debug_module_readdata_from_sa                                  (cpu_linux_jtag_debug_module_readdata_from_sa),
      .d1_cpu_linux_jtag_debug_module_end_xfer                                       (d1_cpu_linux_jtag_debug_module_end_xfer),
      .reset_n                                                                       (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_0 the_Medipix_sopc_burst_0
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_0_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_0_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_0_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_0_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_0_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_0_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_0_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_0_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_0_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_0_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_0_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_0_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_0_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_0_upstream_byteaddress),
      .upstream_byteenable             (Medipix_sopc_burst_0_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_0_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_0_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_0_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_0_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_0_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_0_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_0_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_0_upstream_writedata)
    );

  Medipix_sopc_burst_1_upstream_arbitrator the_Medipix_sopc_burst_1_upstream
    (
      .Medipix_sopc_burst_1_upstream_address                                               (Medipix_sopc_burst_1_upstream_address),
      .Medipix_sopc_burst_1_upstream_burstcount                                            (Medipix_sopc_burst_1_upstream_burstcount),
      .Medipix_sopc_burst_1_upstream_byteaddress                                           (Medipix_sopc_burst_1_upstream_byteaddress),
      .Medipix_sopc_burst_1_upstream_byteenable                                            (Medipix_sopc_burst_1_upstream_byteenable),
      .Medipix_sopc_burst_1_upstream_debugaccess                                           (Medipix_sopc_burst_1_upstream_debugaccess),
      .Medipix_sopc_burst_1_upstream_read                                                  (Medipix_sopc_burst_1_upstream_read),
      .Medipix_sopc_burst_1_upstream_readdata                                              (Medipix_sopc_burst_1_upstream_readdata),
      .Medipix_sopc_burst_1_upstream_readdata_from_sa                                      (Medipix_sopc_burst_1_upstream_readdata_from_sa),
      .Medipix_sopc_burst_1_upstream_readdatavalid                                         (Medipix_sopc_burst_1_upstream_readdatavalid),
      .Medipix_sopc_burst_1_upstream_waitrequest                                           (Medipix_sopc_burst_1_upstream_waitrequest),
      .Medipix_sopc_burst_1_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_1_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_1_upstream_write                                                 (Medipix_sopc_burst_1_upstream_write),
      .Medipix_sopc_burst_1_upstream_writedata                                             (Medipix_sopc_burst_1_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_1_upstream_end_xfer                                           (d1_Medipix_sopc_burst_1_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_1_downstream_arbitrator the_Medipix_sopc_burst_1_downstream
    (
      .Medipix_sopc_burst_1_downstream_address                                       (Medipix_sopc_burst_1_downstream_address),
      .Medipix_sopc_burst_1_downstream_address_to_slave                              (Medipix_sopc_burst_1_downstream_address_to_slave),
      .Medipix_sopc_burst_1_downstream_burstcount                                    (Medipix_sopc_burst_1_downstream_burstcount),
      .Medipix_sopc_burst_1_downstream_byteenable                                    (Medipix_sopc_burst_1_downstream_byteenable),
      .Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module           (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_latency_counter                               (Medipix_sopc_burst_1_downstream_latency_counter),
      .Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module (Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_read                                          (Medipix_sopc_burst_1_downstream_read),
      .Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module   (Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_readdata                                      (Medipix_sopc_burst_1_downstream_readdata),
      .Medipix_sopc_burst_1_downstream_readdatavalid                                 (Medipix_sopc_burst_1_downstream_readdatavalid),
      .Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module          (Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_reset_n                                       (Medipix_sopc_burst_1_downstream_reset_n),
      .Medipix_sopc_burst_1_downstream_waitrequest                                   (Medipix_sopc_burst_1_downstream_waitrequest),
      .Medipix_sopc_burst_1_downstream_write                                         (Medipix_sopc_burst_1_downstream_write),
      .Medipix_sopc_burst_1_downstream_writedata                                     (Medipix_sopc_burst_1_downstream_writedata),
      .clk                                                                           (ram_aux_half_rate_clk_out),
      .cpu_linux_jtag_debug_module_readdata_from_sa                                  (cpu_linux_jtag_debug_module_readdata_from_sa),
      .d1_cpu_linux_jtag_debug_module_end_xfer                                       (d1_cpu_linux_jtag_debug_module_end_xfer),
      .reset_n                                                                       (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_1 the_Medipix_sopc_burst_1
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_1_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_1_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_1_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_1_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_1_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_1_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_1_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_1_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_1_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_1_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_1_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_1_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_1_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_1_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_1_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_1_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_1_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_1_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_1_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_1_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_1_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_1_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_1_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_1_upstream_writedata)
    );

  Medipix_sopc_burst_10_upstream_arbitrator the_Medipix_sopc_burst_10_upstream
    (
      .Medipix_sopc_burst_10_upstream_address                                              (Medipix_sopc_burst_10_upstream_address),
      .Medipix_sopc_burst_10_upstream_burstcount                                           (Medipix_sopc_burst_10_upstream_burstcount),
      .Medipix_sopc_burst_10_upstream_byteaddress                                          (Medipix_sopc_burst_10_upstream_byteaddress),
      .Medipix_sopc_burst_10_upstream_byteenable                                           (Medipix_sopc_burst_10_upstream_byteenable),
      .Medipix_sopc_burst_10_upstream_debugaccess                                          (Medipix_sopc_burst_10_upstream_debugaccess),
      .Medipix_sopc_burst_10_upstream_read                                                 (Medipix_sopc_burst_10_upstream_read),
      .Medipix_sopc_burst_10_upstream_readdata                                             (Medipix_sopc_burst_10_upstream_readdata),
      .Medipix_sopc_burst_10_upstream_readdata_from_sa                                     (Medipix_sopc_burst_10_upstream_readdata_from_sa),
      .Medipix_sopc_burst_10_upstream_readdatavalid                                        (Medipix_sopc_burst_10_upstream_readdatavalid),
      .Medipix_sopc_burst_10_upstream_waitrequest                                          (Medipix_sopc_burst_10_upstream_waitrequest),
      .Medipix_sopc_burst_10_upstream_waitrequest_from_sa                                  (Medipix_sopc_burst_10_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_10_upstream_write                                                (Medipix_sopc_burst_10_upstream_write),
      .Medipix_sopc_burst_10_upstream_writedata                                            (Medipix_sopc_burst_10_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream                        (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream              (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream                (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream                       (cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_10_upstream_end_xfer                                          (d1_Medipix_sopc_burst_10_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_10_downstream_arbitrator the_Medipix_sopc_burst_10_downstream
    (
      .Medipix_sopc_burst_10_downstream_address                                  (Medipix_sopc_burst_10_downstream_address),
      .Medipix_sopc_burst_10_downstream_address_to_slave                         (Medipix_sopc_burst_10_downstream_address_to_slave),
      .Medipix_sopc_burst_10_downstream_burstcount                               (Medipix_sopc_burst_10_downstream_burstcount),
      .Medipix_sopc_burst_10_downstream_byteenable                               (Medipix_sopc_burst_10_downstream_byteenable),
      .Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port           (Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_latency_counter                          (Medipix_sopc_burst_10_downstream_latency_counter),
      .Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port (Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_read                                     (Medipix_sopc_burst_10_downstream_read),
      .Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port   (Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_readdata                                 (Medipix_sopc_burst_10_downstream_readdata),
      .Medipix_sopc_burst_10_downstream_readdatavalid                            (Medipix_sopc_burst_10_downstream_readdatavalid),
      .Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port          (Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_reset_n                                  (Medipix_sopc_burst_10_downstream_reset_n),
      .Medipix_sopc_burst_10_downstream_waitrequest                              (Medipix_sopc_burst_10_downstream_waitrequest),
      .Medipix_sopc_burst_10_downstream_write                                    (Medipix_sopc_burst_10_downstream_write),
      .Medipix_sopc_burst_10_downstream_writedata                                (Medipix_sopc_burst_10_downstream_writedata),
      .clk                                                                       (ram_aux_half_rate_clk_out),
      .d1_spi_0_spi_control_port_end_xfer                                        (d1_spi_0_spi_control_port_end_xfer),
      .reset_n                                                                   (ram_aux_half_rate_clk_out_reset_n),
      .spi_0_spi_control_port_readdata_from_sa                                   (spi_0_spi_control_port_readdata_from_sa)
    );

  Medipix_sopc_burst_10 the_Medipix_sopc_burst_10
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_10_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_10_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_10_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_10_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_10_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_10_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_10_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_10_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_10_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_10_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_10_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_10_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_10_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_10_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_10_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_10_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_10_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_10_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_10_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_10_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_10_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_10_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_10_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_10_upstream_writedata)
    );

  Medipix_sopc_burst_11_upstream_arbitrator the_Medipix_sopc_burst_11_upstream
    (
      .Medipix_sopc_burst_11_upstream_address                                              (Medipix_sopc_burst_11_upstream_address),
      .Medipix_sopc_burst_11_upstream_burstcount                                           (Medipix_sopc_burst_11_upstream_burstcount),
      .Medipix_sopc_burst_11_upstream_byteaddress                                          (Medipix_sopc_burst_11_upstream_byteaddress),
      .Medipix_sopc_burst_11_upstream_byteenable                                           (Medipix_sopc_burst_11_upstream_byteenable),
      .Medipix_sopc_burst_11_upstream_debugaccess                                          (Medipix_sopc_burst_11_upstream_debugaccess),
      .Medipix_sopc_burst_11_upstream_read                                                 (Medipix_sopc_burst_11_upstream_read),
      .Medipix_sopc_burst_11_upstream_readdata                                             (Medipix_sopc_burst_11_upstream_readdata),
      .Medipix_sopc_burst_11_upstream_readdata_from_sa                                     (Medipix_sopc_burst_11_upstream_readdata_from_sa),
      .Medipix_sopc_burst_11_upstream_readdatavalid                                        (Medipix_sopc_burst_11_upstream_readdatavalid),
      .Medipix_sopc_burst_11_upstream_waitrequest                                          (Medipix_sopc_burst_11_upstream_waitrequest),
      .Medipix_sopc_burst_11_upstream_waitrequest_from_sa                                  (Medipix_sopc_burst_11_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_11_upstream_write                                                (Medipix_sopc_burst_11_upstream_write),
      .Medipix_sopc_burst_11_upstream_writedata                                            (Medipix_sopc_burst_11_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream                        (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream              (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream                (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream                       (cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_11_upstream_end_xfer                                          (d1_Medipix_sopc_burst_11_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_11_downstream_arbitrator the_Medipix_sopc_burst_11_downstream
    (
      .Medipix_sopc_burst_11_downstream_address                     (Medipix_sopc_burst_11_downstream_address),
      .Medipix_sopc_burst_11_downstream_address_to_slave            (Medipix_sopc_burst_11_downstream_address_to_slave),
      .Medipix_sopc_burst_11_downstream_burstcount                  (Medipix_sopc_burst_11_downstream_burstcount),
      .Medipix_sopc_burst_11_downstream_byteenable                  (Medipix_sopc_burst_11_downstream_byteenable),
      .Medipix_sopc_burst_11_downstream_granted_uart_0_s1           (Medipix_sopc_burst_11_downstream_granted_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_latency_counter             (Medipix_sopc_burst_11_downstream_latency_counter),
      .Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1 (Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_read                        (Medipix_sopc_burst_11_downstream_read),
      .Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1   (Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_readdata                    (Medipix_sopc_burst_11_downstream_readdata),
      .Medipix_sopc_burst_11_downstream_readdatavalid               (Medipix_sopc_burst_11_downstream_readdatavalid),
      .Medipix_sopc_burst_11_downstream_requests_uart_0_s1          (Medipix_sopc_burst_11_downstream_requests_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_reset_n                     (Medipix_sopc_burst_11_downstream_reset_n),
      .Medipix_sopc_burst_11_downstream_waitrequest                 (Medipix_sopc_burst_11_downstream_waitrequest),
      .Medipix_sopc_burst_11_downstream_write                       (Medipix_sopc_burst_11_downstream_write),
      .Medipix_sopc_burst_11_downstream_writedata                   (Medipix_sopc_burst_11_downstream_writedata),
      .clk                                                          (ram_aux_half_rate_clk_out),
      .d1_uart_0_s1_end_xfer                                        (d1_uart_0_s1_end_xfer),
      .reset_n                                                      (ram_aux_half_rate_clk_out_reset_n),
      .uart_0_s1_readdata_from_sa                                   (uart_0_s1_readdata_from_sa)
    );

  Medipix_sopc_burst_11 the_Medipix_sopc_burst_11
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_11_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_11_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_11_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_11_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_11_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_11_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_11_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_11_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_11_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_11_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_11_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_11_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_11_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_11_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_11_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_11_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_11_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_11_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_11_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_11_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_11_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_11_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_11_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_11_upstream_writedata)
    );

  Medipix_sopc_burst_2_upstream_arbitrator the_Medipix_sopc_burst_2_upstream
    (
      .Medipix_sopc_burst_2_upstream_address                                               (Medipix_sopc_burst_2_upstream_address),
      .Medipix_sopc_burst_2_upstream_burstcount                                            (Medipix_sopc_burst_2_upstream_burstcount),
      .Medipix_sopc_burst_2_upstream_byteaddress                                           (Medipix_sopc_burst_2_upstream_byteaddress),
      .Medipix_sopc_burst_2_upstream_byteenable                                            (Medipix_sopc_burst_2_upstream_byteenable),
      .Medipix_sopc_burst_2_upstream_debugaccess                                           (Medipix_sopc_burst_2_upstream_debugaccess),
      .Medipix_sopc_burst_2_upstream_read                                                  (Medipix_sopc_burst_2_upstream_read),
      .Medipix_sopc_burst_2_upstream_readdata                                              (Medipix_sopc_burst_2_upstream_readdata),
      .Medipix_sopc_burst_2_upstream_readdata_from_sa                                      (Medipix_sopc_burst_2_upstream_readdata_from_sa),
      .Medipix_sopc_burst_2_upstream_readdatavalid                                         (Medipix_sopc_burst_2_upstream_readdatavalid),
      .Medipix_sopc_burst_2_upstream_waitrequest                                           (Medipix_sopc_burst_2_upstream_waitrequest),
      .Medipix_sopc_burst_2_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_2_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_2_upstream_write                                                 (Medipix_sopc_burst_2_upstream_write),
      .Medipix_sopc_burst_2_upstream_writedata                                             (Medipix_sopc_burst_2_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_2_upstream_end_xfer                                           (d1_Medipix_sopc_burst_2_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_2_downstream_arbitrator the_Medipix_sopc_burst_2_downstream
    (
      .Medipix_sopc_burst_2_downstream_address                                         (Medipix_sopc_burst_2_downstream_address),
      .Medipix_sopc_burst_2_downstream_address_to_slave                                (Medipix_sopc_burst_2_downstream_address_to_slave),
      .Medipix_sopc_burst_2_downstream_burstcount                                      (Medipix_sopc_burst_2_downstream_burstcount),
      .Medipix_sopc_burst_2_downstream_byteenable                                      (Medipix_sopc_burst_2_downstream_byteenable),
      .Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave           (Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_latency_counter                                 (Medipix_sopc_burst_2_downstream_latency_counter),
      .Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave (Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_read                                            (Medipix_sopc_burst_2_downstream_read),
      .Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave   (Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_readdata                                        (Medipix_sopc_burst_2_downstream_readdata),
      .Medipix_sopc_burst_2_downstream_readdatavalid                                   (Medipix_sopc_burst_2_downstream_readdatavalid),
      .Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave          (Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_reset_n                                         (Medipix_sopc_burst_2_downstream_reset_n),
      .Medipix_sopc_burst_2_downstream_waitrequest                                     (Medipix_sopc_burst_2_downstream_waitrequest),
      .Medipix_sopc_burst_2_downstream_write                                           (Medipix_sopc_burst_2_downstream_write),
      .Medipix_sopc_burst_2_downstream_writedata                                       (Medipix_sopc_burst_2_downstream_writedata),
      .clk                                                                             (ram_aux_half_rate_clk_out),
      .d1_jtag_uart_0_avalon_jtag_slave_end_xfer                                       (d1_jtag_uart_0_avalon_jtag_slave_end_xfer),
      .jtag_uart_0_avalon_jtag_slave_readdata_from_sa                                  (jtag_uart_0_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa                               (jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa),
      .reset_n                                                                         (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_2 the_Medipix_sopc_burst_2
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_2_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_2_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_2_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_2_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_2_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_2_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_2_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_2_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_2_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_2_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_2_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_2_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_2_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_2_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_2_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_2_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_2_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_2_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_2_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_2_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_2_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_2_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_2_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_2_upstream_writedata)
    );

  Medipix_sopc_burst_3_upstream_arbitrator the_Medipix_sopc_burst_3_upstream
    (
      .Medipix_sopc_burst_3_upstream_address                                               (Medipix_sopc_burst_3_upstream_address),
      .Medipix_sopc_burst_3_upstream_burstcount                                            (Medipix_sopc_burst_3_upstream_burstcount),
      .Medipix_sopc_burst_3_upstream_byteaddress                                           (Medipix_sopc_burst_3_upstream_byteaddress),
      .Medipix_sopc_burst_3_upstream_byteenable                                            (Medipix_sopc_burst_3_upstream_byteenable),
      .Medipix_sopc_burst_3_upstream_debugaccess                                           (Medipix_sopc_burst_3_upstream_debugaccess),
      .Medipix_sopc_burst_3_upstream_read                                                  (Medipix_sopc_burst_3_upstream_read),
      .Medipix_sopc_burst_3_upstream_readdata                                              (Medipix_sopc_burst_3_upstream_readdata),
      .Medipix_sopc_burst_3_upstream_readdata_from_sa                                      (Medipix_sopc_burst_3_upstream_readdata_from_sa),
      .Medipix_sopc_burst_3_upstream_readdatavalid                                         (Medipix_sopc_burst_3_upstream_readdatavalid),
      .Medipix_sopc_burst_3_upstream_waitrequest                                           (Medipix_sopc_burst_3_upstream_waitrequest),
      .Medipix_sopc_burst_3_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_3_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_3_upstream_write                                                 (Medipix_sopc_burst_3_upstream_write),
      .Medipix_sopc_burst_3_upstream_writedata                                             (Medipix_sopc_burst_3_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_3_upstream_end_xfer                                           (d1_Medipix_sopc_burst_3_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_3_downstream_arbitrator the_Medipix_sopc_burst_3_downstream
    (
      .Medipix_sopc_burst_3_downstream_address                           (Medipix_sopc_burst_3_downstream_address),
      .Medipix_sopc_burst_3_downstream_address_to_slave                  (Medipix_sopc_burst_3_downstream_address_to_slave),
      .Medipix_sopc_burst_3_downstream_burstcount                        (Medipix_sopc_burst_3_downstream_burstcount),
      .Medipix_sopc_burst_3_downstream_byteenable                        (Medipix_sopc_burst_3_downstream_byteenable),
      .Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1           (Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_latency_counter                   (Medipix_sopc_burst_3_downstream_latency_counter),
      .Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1 (Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_read                              (Medipix_sopc_burst_3_downstream_read),
      .Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1   (Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_readdata                          (Medipix_sopc_burst_3_downstream_readdata),
      .Medipix_sopc_burst_3_downstream_readdatavalid                     (Medipix_sopc_burst_3_downstream_readdatavalid),
      .Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1          (Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_reset_n                           (Medipix_sopc_burst_3_downstream_reset_n),
      .Medipix_sopc_burst_3_downstream_waitrequest                       (Medipix_sopc_burst_3_downstream_waitrequest),
      .Medipix_sopc_burst_3_downstream_write                             (Medipix_sopc_burst_3_downstream_write),
      .Medipix_sopc_burst_3_downstream_writedata                         (Medipix_sopc_burst_3_downstream_writedata),
      .clk                                                               (ram_aux_half_rate_clk_out),
      .d1_sys_clk_freq_s1_end_xfer                                       (d1_sys_clk_freq_s1_end_xfer),
      .reset_n                                                           (ram_aux_half_rate_clk_out_reset_n),
      .sys_clk_freq_s1_readdata_from_sa                                  (sys_clk_freq_s1_readdata_from_sa)
    );

  Medipix_sopc_burst_3 the_Medipix_sopc_burst_3
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_3_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_3_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_3_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_3_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_3_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_3_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_3_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_3_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_3_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_3_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_3_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_3_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_3_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_3_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_3_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_3_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_3_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_3_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_3_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_3_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_3_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_3_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_3_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_3_upstream_writedata)
    );

  Medipix_sopc_burst_4_upstream_arbitrator the_Medipix_sopc_burst_4_upstream
    (
      .Medipix_sopc_burst_4_upstream_address                                                     (Medipix_sopc_burst_4_upstream_address),
      .Medipix_sopc_burst_4_upstream_byteaddress                                                 (Medipix_sopc_burst_4_upstream_byteaddress),
      .Medipix_sopc_burst_4_upstream_byteenable                                                  (Medipix_sopc_burst_4_upstream_byteenable),
      .Medipix_sopc_burst_4_upstream_debugaccess                                                 (Medipix_sopc_burst_4_upstream_debugaccess),
      .Medipix_sopc_burst_4_upstream_read                                                        (Medipix_sopc_burst_4_upstream_read),
      .Medipix_sopc_burst_4_upstream_readdata                                                    (Medipix_sopc_burst_4_upstream_readdata),
      .Medipix_sopc_burst_4_upstream_readdata_from_sa                                            (Medipix_sopc_burst_4_upstream_readdata_from_sa),
      .Medipix_sopc_burst_4_upstream_readdatavalid                                               (Medipix_sopc_burst_4_upstream_readdatavalid),
      .Medipix_sopc_burst_4_upstream_waitrequest                                                 (Medipix_sopc_burst_4_upstream_waitrequest),
      .Medipix_sopc_burst_4_upstream_waitrequest_from_sa                                         (Medipix_sopc_burst_4_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_4_upstream_write                                                       (Medipix_sopc_burst_4_upstream_write),
      .clk                                                                                       (ram_aux_half_rate_clk_out),
      .cpu_linux_instruction_master_address_to_slave                                             (cpu_linux_instruction_master_address_to_slave),
      .cpu_linux_instruction_master_burstcount                                                   (cpu_linux_instruction_master_burstcount),
      .cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream                        (cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_latency_counter                                              (cpu_linux_instruction_master_latency_counter),
      .cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream              (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_read                                                         (cpu_linux_instruction_master_read),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream                (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register),
      .cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream                       (cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream),
      .d1_Medipix_sopc_burst_4_upstream_end_xfer                                                 (d1_Medipix_sopc_burst_4_upstream_end_xfer),
      .reset_n                                                                                   (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_4_downstream_arbitrator the_Medipix_sopc_burst_4_downstream
    (
      .Medipix_sopc_burst_4_downstream_address                                          (Medipix_sopc_burst_4_downstream_address),
      .Medipix_sopc_burst_4_downstream_address_to_slave                                 (Medipix_sopc_burst_4_downstream_address_to_slave),
      .Medipix_sopc_burst_4_downstream_burstcount                                       (Medipix_sopc_burst_4_downstream_burstcount),
      .Medipix_sopc_burst_4_downstream_byteenable                                       (Medipix_sopc_burst_4_downstream_byteenable),
      .Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1                        (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_latency_counter                                  (Medipix_sopc_burst_4_downstream_latency_counter),
      .Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1              (Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_read                                             (Medipix_sopc_burst_4_downstream_read),
      .Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1                (Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register (Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register),
      .Medipix_sopc_burst_4_downstream_readdata                                         (Medipix_sopc_burst_4_downstream_readdata),
      .Medipix_sopc_burst_4_downstream_readdatavalid                                    (Medipix_sopc_burst_4_downstream_readdatavalid),
      .Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1                       (Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_reset_n                                          (Medipix_sopc_burst_4_downstream_reset_n),
      .Medipix_sopc_burst_4_downstream_waitrequest                                      (Medipix_sopc_burst_4_downstream_waitrequest),
      .Medipix_sopc_burst_4_downstream_write                                            (Medipix_sopc_burst_4_downstream_write),
      .Medipix_sopc_burst_4_downstream_writedata                                        (Medipix_sopc_burst_4_downstream_writedata),
      .clk                                                                              (ram_aux_half_rate_clk_out),
      .clock_crossing_s1_readdata_from_sa                                               (clock_crossing_s1_readdata_from_sa),
      .clock_crossing_s1_waitrequest_from_sa                                            (clock_crossing_s1_waitrequest_from_sa),
      .d1_clock_crossing_s1_end_xfer                                                    (d1_clock_crossing_s1_end_xfer),
      .reset_n                                                                          (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_4 the_Medipix_sopc_burst_4
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_4_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_4_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_4_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_4_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_4_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_4_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_4_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_4_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_4_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_4_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_4_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_4_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_4_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_4_upstream_byteaddress),
      .upstream_byteenable             (Medipix_sopc_burst_4_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_4_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_4_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_4_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_4_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_4_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_4_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_4_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_4_upstream_writedata)
    );

  Medipix_sopc_burst_5_upstream_arbitrator the_Medipix_sopc_burst_5_upstream
    (
      .Medipix_sopc_burst_5_upstream_address                                               (Medipix_sopc_burst_5_upstream_address),
      .Medipix_sopc_burst_5_upstream_burstcount                                            (Medipix_sopc_burst_5_upstream_burstcount),
      .Medipix_sopc_burst_5_upstream_byteaddress                                           (Medipix_sopc_burst_5_upstream_byteaddress),
      .Medipix_sopc_burst_5_upstream_byteenable                                            (Medipix_sopc_burst_5_upstream_byteenable),
      .Medipix_sopc_burst_5_upstream_debugaccess                                           (Medipix_sopc_burst_5_upstream_debugaccess),
      .Medipix_sopc_burst_5_upstream_read                                                  (Medipix_sopc_burst_5_upstream_read),
      .Medipix_sopc_burst_5_upstream_readdata                                              (Medipix_sopc_burst_5_upstream_readdata),
      .Medipix_sopc_burst_5_upstream_readdata_from_sa                                      (Medipix_sopc_burst_5_upstream_readdata_from_sa),
      .Medipix_sopc_burst_5_upstream_readdatavalid                                         (Medipix_sopc_burst_5_upstream_readdatavalid),
      .Medipix_sopc_burst_5_upstream_waitrequest                                           (Medipix_sopc_burst_5_upstream_waitrequest),
      .Medipix_sopc_burst_5_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_5_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_5_upstream_write                                                 (Medipix_sopc_burst_5_upstream_write),
      .Medipix_sopc_burst_5_upstream_writedata                                             (Medipix_sopc_burst_5_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_5_upstream_end_xfer                                           (d1_Medipix_sopc_burst_5_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_5_downstream_arbitrator the_Medipix_sopc_burst_5_downstream
    (
      .Medipix_sopc_burst_5_downstream_address                                          (Medipix_sopc_burst_5_downstream_address),
      .Medipix_sopc_burst_5_downstream_address_to_slave                                 (Medipix_sopc_burst_5_downstream_address_to_slave),
      .Medipix_sopc_burst_5_downstream_burstcount                                       (Medipix_sopc_burst_5_downstream_burstcount),
      .Medipix_sopc_burst_5_downstream_byteenable                                       (Medipix_sopc_burst_5_downstream_byteenable),
      .Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1                        (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_latency_counter                                  (Medipix_sopc_burst_5_downstream_latency_counter),
      .Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1              (Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_read                                             (Medipix_sopc_burst_5_downstream_read),
      .Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1                (Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register (Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register),
      .Medipix_sopc_burst_5_downstream_readdata                                         (Medipix_sopc_burst_5_downstream_readdata),
      .Medipix_sopc_burst_5_downstream_readdatavalid                                    (Medipix_sopc_burst_5_downstream_readdatavalid),
      .Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1                       (Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_reset_n                                          (Medipix_sopc_burst_5_downstream_reset_n),
      .Medipix_sopc_burst_5_downstream_waitrequest                                      (Medipix_sopc_burst_5_downstream_waitrequest),
      .Medipix_sopc_burst_5_downstream_write                                            (Medipix_sopc_burst_5_downstream_write),
      .Medipix_sopc_burst_5_downstream_writedata                                        (Medipix_sopc_burst_5_downstream_writedata),
      .clk                                                                              (ram_aux_half_rate_clk_out),
      .clock_crossing_s1_readdata_from_sa                                               (clock_crossing_s1_readdata_from_sa),
      .clock_crossing_s1_waitrequest_from_sa                                            (clock_crossing_s1_waitrequest_from_sa),
      .d1_clock_crossing_s1_end_xfer                                                    (d1_clock_crossing_s1_end_xfer),
      .reset_n                                                                          (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_5 the_Medipix_sopc_burst_5
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_5_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_5_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_5_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_5_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_5_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_5_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_5_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_5_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_5_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_5_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_5_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_5_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_5_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_5_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_5_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_5_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_5_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_5_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_5_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_5_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_5_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_5_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_5_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_5_upstream_writedata)
    );

  Medipix_sopc_burst_6_upstream_arbitrator the_Medipix_sopc_burst_6_upstream
    (
      .Medipix_sopc_burst_6_upstream_address                                                     (Medipix_sopc_burst_6_upstream_address),
      .Medipix_sopc_burst_6_upstream_byteaddress                                                 (Medipix_sopc_burst_6_upstream_byteaddress),
      .Medipix_sopc_burst_6_upstream_byteenable                                                  (Medipix_sopc_burst_6_upstream_byteenable),
      .Medipix_sopc_burst_6_upstream_debugaccess                                                 (Medipix_sopc_burst_6_upstream_debugaccess),
      .Medipix_sopc_burst_6_upstream_read                                                        (Medipix_sopc_burst_6_upstream_read),
      .Medipix_sopc_burst_6_upstream_readdata                                                    (Medipix_sopc_burst_6_upstream_readdata),
      .Medipix_sopc_burst_6_upstream_readdata_from_sa                                            (Medipix_sopc_burst_6_upstream_readdata_from_sa),
      .Medipix_sopc_burst_6_upstream_readdatavalid                                               (Medipix_sopc_burst_6_upstream_readdatavalid),
      .Medipix_sopc_burst_6_upstream_waitrequest                                                 (Medipix_sopc_burst_6_upstream_waitrequest),
      .Medipix_sopc_burst_6_upstream_waitrequest_from_sa                                         (Medipix_sopc_burst_6_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_6_upstream_write                                                       (Medipix_sopc_burst_6_upstream_write),
      .clk                                                                                       (ram_aux_half_rate_clk_out),
      .cpu_linux_instruction_master_address_to_slave                                             (cpu_linux_instruction_master_address_to_slave),
      .cpu_linux_instruction_master_burstcount                                                   (cpu_linux_instruction_master_burstcount),
      .cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream                        (cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_latency_counter                                              (cpu_linux_instruction_master_latency_counter),
      .cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream              (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_read                                                         (cpu_linux_instruction_master_read),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream                (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register),
      .cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream                       (cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream),
      .d1_Medipix_sopc_burst_6_upstream_end_xfer                                                 (d1_Medipix_sopc_burst_6_upstream_end_xfer),
      .reset_n                                                                                   (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_6_downstream_arbitrator the_Medipix_sopc_burst_6_downstream
    (
      .Medipix_sopc_burst_6_downstream_address                                             (Medipix_sopc_burst_6_downstream_address),
      .Medipix_sopc_burst_6_downstream_address_to_slave                                    (Medipix_sopc_burst_6_downstream_address_to_slave),
      .Medipix_sopc_burst_6_downstream_burstcount                                          (Medipix_sopc_burst_6_downstream_burstcount),
      .Medipix_sopc_burst_6_downstream_byteenable                                          (Medipix_sopc_burst_6_downstream_byteenable),
      .Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port           (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_latency_counter                                     (Medipix_sopc_burst_6_downstream_latency_counter),
      .Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port (Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_read                                                (Medipix_sopc_burst_6_downstream_read),
      .Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port   (Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_readdata                                            (Medipix_sopc_burst_6_downstream_readdata),
      .Medipix_sopc_burst_6_downstream_readdatavalid                                       (Medipix_sopc_burst_6_downstream_readdatavalid),
      .Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port          (Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_reset_n                                             (Medipix_sopc_burst_6_downstream_reset_n),
      .Medipix_sopc_burst_6_downstream_waitrequest                                         (Medipix_sopc_burst_6_downstream_waitrequest),
      .Medipix_sopc_burst_6_downstream_write                                               (Medipix_sopc_burst_6_downstream_write),
      .Medipix_sopc_burst_6_downstream_writedata                                           (Medipix_sopc_burst_6_downstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .d1_epcs_controller_epcs_control_port_end_xfer                                       (d1_epcs_controller_epcs_control_port_end_xfer),
      .epcs_controller_epcs_control_port_readdata_from_sa                                  (epcs_controller_epcs_control_port_readdata_from_sa),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_6 the_Medipix_sopc_burst_6
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_6_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_6_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_6_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_6_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_6_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_6_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_6_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_6_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_6_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_6_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_6_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_6_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_6_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_6_upstream_byteaddress),
      .upstream_byteenable             (Medipix_sopc_burst_6_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_6_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_6_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_6_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_6_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_6_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_6_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_6_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_6_upstream_writedata)
    );

  Medipix_sopc_burst_7_upstream_arbitrator the_Medipix_sopc_burst_7_upstream
    (
      .Medipix_sopc_burst_7_upstream_address                                               (Medipix_sopc_burst_7_upstream_address),
      .Medipix_sopc_burst_7_upstream_burstcount                                            (Medipix_sopc_burst_7_upstream_burstcount),
      .Medipix_sopc_burst_7_upstream_byteaddress                                           (Medipix_sopc_burst_7_upstream_byteaddress),
      .Medipix_sopc_burst_7_upstream_byteenable                                            (Medipix_sopc_burst_7_upstream_byteenable),
      .Medipix_sopc_burst_7_upstream_debugaccess                                           (Medipix_sopc_burst_7_upstream_debugaccess),
      .Medipix_sopc_burst_7_upstream_read                                                  (Medipix_sopc_burst_7_upstream_read),
      .Medipix_sopc_burst_7_upstream_readdata                                              (Medipix_sopc_burst_7_upstream_readdata),
      .Medipix_sopc_burst_7_upstream_readdata_from_sa                                      (Medipix_sopc_burst_7_upstream_readdata_from_sa),
      .Medipix_sopc_burst_7_upstream_readdatavalid                                         (Medipix_sopc_burst_7_upstream_readdatavalid),
      .Medipix_sopc_burst_7_upstream_waitrequest                                           (Medipix_sopc_burst_7_upstream_waitrequest),
      .Medipix_sopc_burst_7_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_7_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_7_upstream_write                                                 (Medipix_sopc_burst_7_upstream_write),
      .Medipix_sopc_burst_7_upstream_writedata                                             (Medipix_sopc_burst_7_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_7_upstream_end_xfer                                           (d1_Medipix_sopc_burst_7_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_7_downstream_arbitrator the_Medipix_sopc_burst_7_downstream
    (
      .Medipix_sopc_burst_7_downstream_address                                             (Medipix_sopc_burst_7_downstream_address),
      .Medipix_sopc_burst_7_downstream_address_to_slave                                    (Medipix_sopc_burst_7_downstream_address_to_slave),
      .Medipix_sopc_burst_7_downstream_burstcount                                          (Medipix_sopc_burst_7_downstream_burstcount),
      .Medipix_sopc_burst_7_downstream_byteenable                                          (Medipix_sopc_burst_7_downstream_byteenable),
      .Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port           (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_latency_counter                                     (Medipix_sopc_burst_7_downstream_latency_counter),
      .Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port (Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_read                                                (Medipix_sopc_burst_7_downstream_read),
      .Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port   (Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_readdata                                            (Medipix_sopc_burst_7_downstream_readdata),
      .Medipix_sopc_burst_7_downstream_readdatavalid                                       (Medipix_sopc_burst_7_downstream_readdatavalid),
      .Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port          (Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_reset_n                                             (Medipix_sopc_burst_7_downstream_reset_n),
      .Medipix_sopc_burst_7_downstream_waitrequest                                         (Medipix_sopc_burst_7_downstream_waitrequest),
      .Medipix_sopc_burst_7_downstream_write                                               (Medipix_sopc_burst_7_downstream_write),
      .Medipix_sopc_burst_7_downstream_writedata                                           (Medipix_sopc_burst_7_downstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .d1_epcs_controller_epcs_control_port_end_xfer                                       (d1_epcs_controller_epcs_control_port_end_xfer),
      .epcs_controller_epcs_control_port_readdata_from_sa                                  (epcs_controller_epcs_control_port_readdata_from_sa),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_7 the_Medipix_sopc_burst_7
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_7_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_7_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_7_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_7_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_7_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_7_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_7_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_7_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_7_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_7_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_7_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_7_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_7_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_7_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_7_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_7_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_7_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_7_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_7_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_7_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_7_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_7_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_7_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_7_upstream_writedata)
    );

  Medipix_sopc_burst_8_upstream_arbitrator the_Medipix_sopc_burst_8_upstream
    (
      .Medipix_sopc_burst_8_upstream_address                                               (Medipix_sopc_burst_8_upstream_address),
      .Medipix_sopc_burst_8_upstream_burstcount                                            (Medipix_sopc_burst_8_upstream_burstcount),
      .Medipix_sopc_burst_8_upstream_byteaddress                                           (Medipix_sopc_burst_8_upstream_byteaddress),
      .Medipix_sopc_burst_8_upstream_byteenable                                            (Medipix_sopc_burst_8_upstream_byteenable),
      .Medipix_sopc_burst_8_upstream_debugaccess                                           (Medipix_sopc_burst_8_upstream_debugaccess),
      .Medipix_sopc_burst_8_upstream_read                                                  (Medipix_sopc_burst_8_upstream_read),
      .Medipix_sopc_burst_8_upstream_readdata                                              (Medipix_sopc_burst_8_upstream_readdata),
      .Medipix_sopc_burst_8_upstream_readdata_from_sa                                      (Medipix_sopc_burst_8_upstream_readdata_from_sa),
      .Medipix_sopc_burst_8_upstream_readdatavalid                                         (Medipix_sopc_burst_8_upstream_readdatavalid),
      .Medipix_sopc_burst_8_upstream_waitrequest                                           (Medipix_sopc_burst_8_upstream_waitrequest),
      .Medipix_sopc_burst_8_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_8_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_8_upstream_write                                                 (Medipix_sopc_burst_8_upstream_write),
      .Medipix_sopc_burst_8_upstream_writedata                                             (Medipix_sopc_burst_8_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_8_upstream_end_xfer                                           (d1_Medipix_sopc_burst_8_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_8_downstream_arbitrator the_Medipix_sopc_burst_8_downstream
    (
      .Medipix_sopc_burst_8_downstream_address                                 (Medipix_sopc_burst_8_downstream_address),
      .Medipix_sopc_burst_8_downstream_address_to_slave                        (Medipix_sopc_burst_8_downstream_address_to_slave),
      .Medipix_sopc_burst_8_downstream_burstcount                              (Medipix_sopc_burst_8_downstream_burstcount),
      .Medipix_sopc_burst_8_downstream_byteenable                              (Medipix_sopc_burst_8_downstream_byteenable),
      .Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port           (Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_latency_counter                         (Medipix_sopc_burst_8_downstream_latency_counter),
      .Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port (Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_read                                    (Medipix_sopc_burst_8_downstream_read),
      .Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port   (Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_readdata                                (Medipix_sopc_burst_8_downstream_readdata),
      .Medipix_sopc_burst_8_downstream_readdatavalid                           (Medipix_sopc_burst_8_downstream_readdatavalid),
      .Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port          (Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_reset_n                                 (Medipix_sopc_burst_8_downstream_reset_n),
      .Medipix_sopc_burst_8_downstream_waitrequest                             (Medipix_sopc_burst_8_downstream_waitrequest),
      .Medipix_sopc_burst_8_downstream_write                                   (Medipix_sopc_burst_8_downstream_write),
      .Medipix_sopc_burst_8_downstream_writedata                               (Medipix_sopc_burst_8_downstream_writedata),
      .clk                                                                     (ram_aux_half_rate_clk_out),
      .d1_igor_mac_control_port_end_xfer                                       (d1_igor_mac_control_port_end_xfer),
      .igor_mac_control_port_readdata_from_sa                                  (igor_mac_control_port_readdata_from_sa),
      .igor_mac_control_port_waitrequest_n_from_sa                             (igor_mac_control_port_waitrequest_n_from_sa),
      .reset_n                                                                 (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_8 the_Medipix_sopc_burst_8
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_8_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_8_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_8_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_8_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_8_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_8_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_8_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_8_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_8_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_8_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_8_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_8_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_8_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_8_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_8_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_8_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_8_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_8_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_8_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_8_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_8_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_8_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_8_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_8_upstream_writedata)
    );

  Medipix_sopc_burst_9_upstream_arbitrator the_Medipix_sopc_burst_9_upstream
    (
      .Medipix_sopc_burst_9_upstream_address                                               (Medipix_sopc_burst_9_upstream_address),
      .Medipix_sopc_burst_9_upstream_burstcount                                            (Medipix_sopc_burst_9_upstream_burstcount),
      .Medipix_sopc_burst_9_upstream_byteaddress                                           (Medipix_sopc_burst_9_upstream_byteaddress),
      .Medipix_sopc_burst_9_upstream_byteenable                                            (Medipix_sopc_burst_9_upstream_byteenable),
      .Medipix_sopc_burst_9_upstream_debugaccess                                           (Medipix_sopc_burst_9_upstream_debugaccess),
      .Medipix_sopc_burst_9_upstream_read                                                  (Medipix_sopc_burst_9_upstream_read),
      .Medipix_sopc_burst_9_upstream_readdata                                              (Medipix_sopc_burst_9_upstream_readdata),
      .Medipix_sopc_burst_9_upstream_readdata_from_sa                                      (Medipix_sopc_burst_9_upstream_readdata_from_sa),
      .Medipix_sopc_burst_9_upstream_readdatavalid                                         (Medipix_sopc_burst_9_upstream_readdatavalid),
      .Medipix_sopc_burst_9_upstream_waitrequest                                           (Medipix_sopc_burst_9_upstream_waitrequest),
      .Medipix_sopc_burst_9_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_9_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_9_upstream_write                                                 (Medipix_sopc_burst_9_upstream_write),
      .Medipix_sopc_burst_9_upstream_writedata                                             (Medipix_sopc_burst_9_upstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_debugaccess                                                   (cpu_linux_data_master_debugaccess),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_9_upstream_end_xfer                                           (d1_Medipix_sopc_burst_9_upstream_end_xfer),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  Medipix_sopc_burst_9_downstream_arbitrator the_Medipix_sopc_burst_9_downstream
    (
      .Medipix_sopc_burst_9_downstream_address                                   (Medipix_sopc_burst_9_downstream_address),
      .Medipix_sopc_burst_9_downstream_address_to_slave                          (Medipix_sopc_burst_9_downstream_address_to_slave),
      .Medipix_sopc_burst_9_downstream_burstcount                                (Medipix_sopc_burst_9_downstream_burstcount),
      .Medipix_sopc_burst_9_downstream_byteenable                                (Medipix_sopc_burst_9_downstream_byteenable),
      .Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0           (Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_latency_counter                           (Medipix_sopc_burst_9_downstream_latency_counter),
      .Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0 (Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_read                                      (Medipix_sopc_burst_9_downstream_read),
      .Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0   (Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_readdata                                  (Medipix_sopc_burst_9_downstream_readdata),
      .Medipix_sopc_burst_9_downstream_readdatavalid                             (Medipix_sopc_burst_9_downstream_readdatavalid),
      .Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0          (Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_reset_n                                   (Medipix_sopc_burst_9_downstream_reset_n),
      .Medipix_sopc_burst_9_downstream_waitrequest                               (Medipix_sopc_burst_9_downstream_waitrequest),
      .Medipix_sopc_burst_9_downstream_write                                     (Medipix_sopc_burst_9_downstream_write),
      .Medipix_sopc_burst_9_downstream_writedata                                 (Medipix_sopc_burst_9_downstream_writedata),
      .clk                                                                       (ram_aux_half_rate_clk_out),
      .d1_tx_table_avalon_slave_0_end_xfer                                       (d1_tx_table_avalon_slave_0_end_xfer),
      .reset_n                                                                   (ram_aux_half_rate_clk_out_reset_n),
      .tx_table_avalon_slave_0_readdata_from_sa                                  (tx_table_avalon_slave_0_readdata_from_sa)
    );

  Medipix_sopc_burst_9 the_Medipix_sopc_burst_9
    (
      .clk                             (ram_aux_half_rate_clk_out),
      .downstream_readdata             (Medipix_sopc_burst_9_downstream_readdata),
      .downstream_readdatavalid        (Medipix_sopc_burst_9_downstream_readdatavalid),
      .downstream_waitrequest          (Medipix_sopc_burst_9_downstream_waitrequest),
      .reg_downstream_address          (Medipix_sopc_burst_9_downstream_address),
      .reg_downstream_arbitrationshare (Medipix_sopc_burst_9_downstream_arbitrationshare),
      .reg_downstream_burstcount       (Medipix_sopc_burst_9_downstream_burstcount),
      .reg_downstream_byteenable       (Medipix_sopc_burst_9_downstream_byteenable),
      .reg_downstream_debugaccess      (Medipix_sopc_burst_9_downstream_debugaccess),
      .reg_downstream_nativeaddress    (Medipix_sopc_burst_9_downstream_nativeaddress),
      .reg_downstream_read             (Medipix_sopc_burst_9_downstream_read),
      .reg_downstream_write            (Medipix_sopc_burst_9_downstream_write),
      .reg_downstream_writedata        (Medipix_sopc_burst_9_downstream_writedata),
      .reset_n                         (Medipix_sopc_burst_9_downstream_reset_n),
      .upstream_address                (Medipix_sopc_burst_9_upstream_byteaddress),
      .upstream_burstcount             (Medipix_sopc_burst_9_upstream_burstcount),
      .upstream_byteenable             (Medipix_sopc_burst_9_upstream_byteenable),
      .upstream_debugaccess            (Medipix_sopc_burst_9_upstream_debugaccess),
      .upstream_nativeaddress          (Medipix_sopc_burst_9_upstream_address),
      .upstream_read                   (Medipix_sopc_burst_9_upstream_read),
      .upstream_readdata               (Medipix_sopc_burst_9_upstream_readdata),
      .upstream_readdatavalid          (Medipix_sopc_burst_9_upstream_readdatavalid),
      .upstream_waitrequest            (Medipix_sopc_burst_9_upstream_waitrequest),
      .upstream_write                  (Medipix_sopc_burst_9_upstream_write),
      .upstream_writedata              (Medipix_sopc_burst_9_upstream_writedata)
    );

  clock_crossing_s1_arbitrator the_clock_crossing_s1
    (
      .Medipix_sopc_burst_4_downstream_address_to_slave                                 (Medipix_sopc_burst_4_downstream_address_to_slave),
      .Medipix_sopc_burst_4_downstream_arbitrationshare                                 (Medipix_sopc_burst_4_downstream_arbitrationshare),
      .Medipix_sopc_burst_4_downstream_burstcount                                       (Medipix_sopc_burst_4_downstream_burstcount),
      .Medipix_sopc_burst_4_downstream_byteenable                                       (Medipix_sopc_burst_4_downstream_byteenable),
      .Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1                        (Medipix_sopc_burst_4_downstream_granted_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_latency_counter                                  (Medipix_sopc_burst_4_downstream_latency_counter),
      .Medipix_sopc_burst_4_downstream_nativeaddress                                    (Medipix_sopc_burst_4_downstream_nativeaddress),
      .Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1              (Medipix_sopc_burst_4_downstream_qualified_request_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_read                                             (Medipix_sopc_burst_4_downstream_read),
      .Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1                (Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register (Medipix_sopc_burst_4_downstream_read_data_valid_clock_crossing_s1_shift_register),
      .Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1                       (Medipix_sopc_burst_4_downstream_requests_clock_crossing_s1),
      .Medipix_sopc_burst_4_downstream_write                                            (Medipix_sopc_burst_4_downstream_write),
      .Medipix_sopc_burst_4_downstream_writedata                                        (Medipix_sopc_burst_4_downstream_writedata),
      .Medipix_sopc_burst_5_downstream_address_to_slave                                 (Medipix_sopc_burst_5_downstream_address_to_slave),
      .Medipix_sopc_burst_5_downstream_arbitrationshare                                 (Medipix_sopc_burst_5_downstream_arbitrationshare),
      .Medipix_sopc_burst_5_downstream_burstcount                                       (Medipix_sopc_burst_5_downstream_burstcount),
      .Medipix_sopc_burst_5_downstream_byteenable                                       (Medipix_sopc_burst_5_downstream_byteenable),
      .Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1                        (Medipix_sopc_burst_5_downstream_granted_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_latency_counter                                  (Medipix_sopc_burst_5_downstream_latency_counter),
      .Medipix_sopc_burst_5_downstream_nativeaddress                                    (Medipix_sopc_burst_5_downstream_nativeaddress),
      .Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1              (Medipix_sopc_burst_5_downstream_qualified_request_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_read                                             (Medipix_sopc_burst_5_downstream_read),
      .Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1                (Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register (Medipix_sopc_burst_5_downstream_read_data_valid_clock_crossing_s1_shift_register),
      .Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1                       (Medipix_sopc_burst_5_downstream_requests_clock_crossing_s1),
      .Medipix_sopc_burst_5_downstream_write                                            (Medipix_sopc_burst_5_downstream_write),
      .Medipix_sopc_burst_5_downstream_writedata                                        (Medipix_sopc_burst_5_downstream_writedata),
      .clk                                                                              (ram_aux_half_rate_clk_out),
      .clock_crossing_s1_address                                                        (clock_crossing_s1_address),
      .clock_crossing_s1_byteenable                                                     (clock_crossing_s1_byteenable),
      .clock_crossing_s1_endofpacket                                                    (clock_crossing_s1_endofpacket),
      .clock_crossing_s1_endofpacket_from_sa                                            (clock_crossing_s1_endofpacket_from_sa),
      .clock_crossing_s1_nativeaddress                                                  (clock_crossing_s1_nativeaddress),
      .clock_crossing_s1_read                                                           (clock_crossing_s1_read),
      .clock_crossing_s1_readdata                                                       (clock_crossing_s1_readdata),
      .clock_crossing_s1_readdata_from_sa                                               (clock_crossing_s1_readdata_from_sa),
      .clock_crossing_s1_readdatavalid                                                  (clock_crossing_s1_readdatavalid),
      .clock_crossing_s1_reset_n                                                        (clock_crossing_s1_reset_n),
      .clock_crossing_s1_waitrequest                                                    (clock_crossing_s1_waitrequest),
      .clock_crossing_s1_waitrequest_from_sa                                            (clock_crossing_s1_waitrequest_from_sa),
      .clock_crossing_s1_write                                                          (clock_crossing_s1_write),
      .clock_crossing_s1_writedata                                                      (clock_crossing_s1_writedata),
      .d1_clock_crossing_s1_end_xfer                                                    (d1_clock_crossing_s1_end_xfer),
      .igor_mac_rx_master_address_to_slave                                              (igor_mac_rx_master_address_to_slave),
      .igor_mac_rx_master_byteenable                                                    (igor_mac_rx_master_byteenable),
      .igor_mac_rx_master_granted_clock_crossing_s1                                     (igor_mac_rx_master_granted_clock_crossing_s1),
      .igor_mac_rx_master_qualified_request_clock_crossing_s1                           (igor_mac_rx_master_qualified_request_clock_crossing_s1),
      .igor_mac_rx_master_requests_clock_crossing_s1                                    (igor_mac_rx_master_requests_clock_crossing_s1),
      .igor_mac_rx_master_write                                                         (igor_mac_rx_master_write),
      .igor_mac_rx_master_writedata                                                     (igor_mac_rx_master_writedata),
      .igor_mac_tx_master_address_to_slave                                              (igor_mac_tx_master_address_to_slave),
      .igor_mac_tx_master_granted_clock_crossing_s1                                     (igor_mac_tx_master_granted_clock_crossing_s1),
      .igor_mac_tx_master_latency_counter                                               (igor_mac_tx_master_latency_counter),
      .igor_mac_tx_master_qualified_request_clock_crossing_s1                           (igor_mac_tx_master_qualified_request_clock_crossing_s1),
      .igor_mac_tx_master_read                                                          (igor_mac_tx_master_read),
      .igor_mac_tx_master_read_data_valid_clock_crossing_s1                             (igor_mac_tx_master_read_data_valid_clock_crossing_s1),
      .igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register              (igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register),
      .igor_mac_tx_master_requests_clock_crossing_s1                                    (igor_mac_tx_master_requests_clock_crossing_s1),
      .reset_n                                                                          (ram_aux_half_rate_clk_out_reset_n)
    );

  clock_crossing_m1_arbitrator the_clock_crossing_m1
    (
      .clk                                                     (ram_phy_clk_out),
      .clock_crossing_m1_address                               (clock_crossing_m1_address),
      .clock_crossing_m1_address_to_slave                      (clock_crossing_m1_address_to_slave),
      .clock_crossing_m1_byteenable                            (clock_crossing_m1_byteenable),
      .clock_crossing_m1_granted_ram_s1                        (clock_crossing_m1_granted_ram_s1),
      .clock_crossing_m1_latency_counter                       (clock_crossing_m1_latency_counter),
      .clock_crossing_m1_qualified_request_ram_s1              (clock_crossing_m1_qualified_request_ram_s1),
      .clock_crossing_m1_read                                  (clock_crossing_m1_read),
      .clock_crossing_m1_read_data_valid_ram_s1                (clock_crossing_m1_read_data_valid_ram_s1),
      .clock_crossing_m1_read_data_valid_ram_s1_shift_register (clock_crossing_m1_read_data_valid_ram_s1_shift_register),
      .clock_crossing_m1_readdata                              (clock_crossing_m1_readdata),
      .clock_crossing_m1_readdatavalid                         (clock_crossing_m1_readdatavalid),
      .clock_crossing_m1_requests_ram_s1                       (clock_crossing_m1_requests_ram_s1),
      .clock_crossing_m1_reset_n                               (clock_crossing_m1_reset_n),
      .clock_crossing_m1_waitrequest                           (clock_crossing_m1_waitrequest),
      .clock_crossing_m1_write                                 (clock_crossing_m1_write),
      .clock_crossing_m1_writedata                             (clock_crossing_m1_writedata),
      .d1_ram_s1_end_xfer                                      (d1_ram_s1_end_xfer),
      .ram_s1_readdata_from_sa                                 (ram_s1_readdata_from_sa),
      .ram_s1_waitrequest_n_from_sa                            (ram_s1_waitrequest_n_from_sa),
      .reset_n                                                 (ram_phy_clk_out_reset_n)
    );

  clock_crossing the_clock_crossing
    (
      .master_address       (clock_crossing_m1_address),
      .master_byteenable    (clock_crossing_m1_byteenable),
      .master_clk           (ram_phy_clk_out),
      .master_endofpacket   (clock_crossing_m1_endofpacket),
      .master_nativeaddress (clock_crossing_m1_nativeaddress),
      .master_read          (clock_crossing_m1_read),
      .master_readdata      (clock_crossing_m1_readdata),
      .master_readdatavalid (clock_crossing_m1_readdatavalid),
      .master_reset_n       (clock_crossing_m1_reset_n),
      .master_waitrequest   (clock_crossing_m1_waitrequest),
      .master_write         (clock_crossing_m1_write),
      .master_writedata     (clock_crossing_m1_writedata),
      .slave_address        (clock_crossing_s1_address),
      .slave_byteenable     (clock_crossing_s1_byteenable),
      .slave_clk            (ram_aux_half_rate_clk_out),
      .slave_endofpacket    (clock_crossing_s1_endofpacket),
      .slave_nativeaddress  (clock_crossing_s1_nativeaddress),
      .slave_read           (clock_crossing_s1_read),
      .slave_readdata       (clock_crossing_s1_readdata),
      .slave_readdatavalid  (clock_crossing_s1_readdatavalid),
      .slave_reset_n        (clock_crossing_s1_reset_n),
      .slave_waitrequest    (clock_crossing_s1_waitrequest),
      .slave_write          (clock_crossing_s1_write),
      .slave_writedata      (clock_crossing_s1_writedata)
    );

  cpu_linux_jtag_debug_module_arbitrator the_cpu_linux_jtag_debug_module
    (
      .Medipix_sopc_burst_0_downstream_address_to_slave                              (Medipix_sopc_burst_0_downstream_address_to_slave),
      .Medipix_sopc_burst_0_downstream_arbitrationshare                              (Medipix_sopc_burst_0_downstream_arbitrationshare),
      .Medipix_sopc_burst_0_downstream_burstcount                                    (Medipix_sopc_burst_0_downstream_burstcount),
      .Medipix_sopc_burst_0_downstream_byteenable                                    (Medipix_sopc_burst_0_downstream_byteenable),
      .Medipix_sopc_burst_0_downstream_debugaccess                                   (Medipix_sopc_burst_0_downstream_debugaccess),
      .Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module           (Medipix_sopc_burst_0_downstream_granted_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_latency_counter                               (Medipix_sopc_burst_0_downstream_latency_counter),
      .Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module (Medipix_sopc_burst_0_downstream_qualified_request_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_read                                          (Medipix_sopc_burst_0_downstream_read),
      .Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module   (Medipix_sopc_burst_0_downstream_read_data_valid_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module          (Medipix_sopc_burst_0_downstream_requests_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_0_downstream_write                                         (Medipix_sopc_burst_0_downstream_write),
      .Medipix_sopc_burst_0_downstream_writedata                                     (Medipix_sopc_burst_0_downstream_writedata),
      .Medipix_sopc_burst_1_downstream_address_to_slave                              (Medipix_sopc_burst_1_downstream_address_to_slave),
      .Medipix_sopc_burst_1_downstream_arbitrationshare                              (Medipix_sopc_burst_1_downstream_arbitrationshare),
      .Medipix_sopc_burst_1_downstream_burstcount                                    (Medipix_sopc_burst_1_downstream_burstcount),
      .Medipix_sopc_burst_1_downstream_byteenable                                    (Medipix_sopc_burst_1_downstream_byteenable),
      .Medipix_sopc_burst_1_downstream_debugaccess                                   (Medipix_sopc_burst_1_downstream_debugaccess),
      .Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module           (Medipix_sopc_burst_1_downstream_granted_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_latency_counter                               (Medipix_sopc_burst_1_downstream_latency_counter),
      .Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module (Medipix_sopc_burst_1_downstream_qualified_request_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_read                                          (Medipix_sopc_burst_1_downstream_read),
      .Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module   (Medipix_sopc_burst_1_downstream_read_data_valid_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module          (Medipix_sopc_burst_1_downstream_requests_cpu_linux_jtag_debug_module),
      .Medipix_sopc_burst_1_downstream_write                                         (Medipix_sopc_burst_1_downstream_write),
      .Medipix_sopc_burst_1_downstream_writedata                                     (Medipix_sopc_burst_1_downstream_writedata),
      .clk                                                                           (ram_aux_half_rate_clk_out),
      .cpu_linux_jtag_debug_module_address                                           (cpu_linux_jtag_debug_module_address),
      .cpu_linux_jtag_debug_module_begintransfer                                     (cpu_linux_jtag_debug_module_begintransfer),
      .cpu_linux_jtag_debug_module_byteenable                                        (cpu_linux_jtag_debug_module_byteenable),
      .cpu_linux_jtag_debug_module_chipselect                                        (cpu_linux_jtag_debug_module_chipselect),
      .cpu_linux_jtag_debug_module_debugaccess                                       (cpu_linux_jtag_debug_module_debugaccess),
      .cpu_linux_jtag_debug_module_readdata                                          (cpu_linux_jtag_debug_module_readdata),
      .cpu_linux_jtag_debug_module_readdata_from_sa                                  (cpu_linux_jtag_debug_module_readdata_from_sa),
      .cpu_linux_jtag_debug_module_reset_n                                           (cpu_linux_jtag_debug_module_reset_n),
      .cpu_linux_jtag_debug_module_resetrequest                                      (cpu_linux_jtag_debug_module_resetrequest),
      .cpu_linux_jtag_debug_module_resetrequest_from_sa                              (cpu_linux_jtag_debug_module_resetrequest_from_sa),
      .cpu_linux_jtag_debug_module_write                                             (cpu_linux_jtag_debug_module_write),
      .cpu_linux_jtag_debug_module_writedata                                         (cpu_linux_jtag_debug_module_writedata),
      .d1_cpu_linux_jtag_debug_module_end_xfer                                       (d1_cpu_linux_jtag_debug_module_end_xfer),
      .reset_n                                                                       (ram_aux_half_rate_clk_out_reset_n)
    );

  cpu_linux_data_master_arbitrator the_cpu_linux_data_master
    (
      .Medipix_sopc_burst_10_upstream_readdata_from_sa                                     (Medipix_sopc_burst_10_upstream_readdata_from_sa),
      .Medipix_sopc_burst_10_upstream_waitrequest_from_sa                                  (Medipix_sopc_burst_10_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_11_upstream_readdata_from_sa                                     (Medipix_sopc_burst_11_upstream_readdata_from_sa),
      .Medipix_sopc_burst_11_upstream_waitrequest_from_sa                                  (Medipix_sopc_burst_11_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_1_upstream_readdata_from_sa                                      (Medipix_sopc_burst_1_upstream_readdata_from_sa),
      .Medipix_sopc_burst_1_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_1_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_2_upstream_readdata_from_sa                                      (Medipix_sopc_burst_2_upstream_readdata_from_sa),
      .Medipix_sopc_burst_2_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_2_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_3_upstream_readdata_from_sa                                      (Medipix_sopc_burst_3_upstream_readdata_from_sa),
      .Medipix_sopc_burst_3_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_3_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_5_upstream_readdata_from_sa                                      (Medipix_sopc_burst_5_upstream_readdata_from_sa),
      .Medipix_sopc_burst_5_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_5_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_7_upstream_readdata_from_sa                                      (Medipix_sopc_burst_7_upstream_readdata_from_sa),
      .Medipix_sopc_burst_7_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_7_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_8_upstream_readdata_from_sa                                      (Medipix_sopc_burst_8_upstream_readdata_from_sa),
      .Medipix_sopc_burst_8_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_8_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_9_upstream_readdata_from_sa                                      (Medipix_sopc_burst_9_upstream_readdata_from_sa),
      .Medipix_sopc_burst_9_upstream_waitrequest_from_sa                                   (Medipix_sopc_burst_9_upstream_waitrequest_from_sa),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .cpu_linux_data_master_address                                                       (cpu_linux_data_master_address),
      .cpu_linux_data_master_address_to_slave                                              (cpu_linux_data_master_address_to_slave),
      .cpu_linux_data_master_burstcount                                                    (cpu_linux_data_master_burstcount),
      .cpu_linux_data_master_byteenable                                                    (cpu_linux_data_master_byteenable),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream                        (cpu_linux_data_master_granted_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream                        (cpu_linux_data_master_granted_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream                         (cpu_linux_data_master_granted_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_irq                                                           (cpu_linux_data_master_irq),
      .cpu_linux_data_master_latency_counter                                               (cpu_linux_data_master_latency_counter),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream              (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream              (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream               (cpu_linux_data_master_qualified_request_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_read                                                          (cpu_linux_data_master_read),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream                (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_10_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream                (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_11_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_1_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_2_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_3_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_5_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_7_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_8_upstream_shift_register),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream                 (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register  (cpu_linux_data_master_read_data_valid_Medipix_sopc_burst_9_upstream_shift_register),
      .cpu_linux_data_master_readdata                                                      (cpu_linux_data_master_readdata),
      .cpu_linux_data_master_readdatavalid                                                 (cpu_linux_data_master_readdatavalid),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream                       (cpu_linux_data_master_requests_Medipix_sopc_burst_10_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream                       (cpu_linux_data_master_requests_Medipix_sopc_burst_11_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_1_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_2_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_3_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_5_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_7_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_8_upstream),
      .cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream                        (cpu_linux_data_master_requests_Medipix_sopc_burst_9_upstream),
      .cpu_linux_data_master_waitrequest                                                   (cpu_linux_data_master_waitrequest),
      .cpu_linux_data_master_write                                                         (cpu_linux_data_master_write),
      .cpu_linux_data_master_writedata                                                     (cpu_linux_data_master_writedata),
      .d1_Medipix_sopc_burst_10_upstream_end_xfer                                          (d1_Medipix_sopc_burst_10_upstream_end_xfer),
      .d1_Medipix_sopc_burst_11_upstream_end_xfer                                          (d1_Medipix_sopc_burst_11_upstream_end_xfer),
      .d1_Medipix_sopc_burst_1_upstream_end_xfer                                           (d1_Medipix_sopc_burst_1_upstream_end_xfer),
      .d1_Medipix_sopc_burst_2_upstream_end_xfer                                           (d1_Medipix_sopc_burst_2_upstream_end_xfer),
      .d1_Medipix_sopc_burst_3_upstream_end_xfer                                           (d1_Medipix_sopc_burst_3_upstream_end_xfer),
      .d1_Medipix_sopc_burst_5_upstream_end_xfer                                           (d1_Medipix_sopc_burst_5_upstream_end_xfer),
      .d1_Medipix_sopc_burst_7_upstream_end_xfer                                           (d1_Medipix_sopc_burst_7_upstream_end_xfer),
      .d1_Medipix_sopc_burst_8_upstream_end_xfer                                           (d1_Medipix_sopc_burst_8_upstream_end_xfer),
      .d1_Medipix_sopc_burst_9_upstream_end_xfer                                           (d1_Medipix_sopc_burst_9_upstream_end_xfer),
      .epcs_controller_epcs_control_port_irq_from_sa                                       (epcs_controller_epcs_control_port_irq_from_sa),
      .igor_mac_control_port_irq_from_sa                                                   (igor_mac_control_port_irq_from_sa),
      .jtag_uart_0_avalon_jtag_slave_irq_from_sa                                           (jtag_uart_0_avalon_jtag_slave_irq_from_sa),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n),
      .spi_0_spi_control_port_irq_from_sa                                                  (spi_0_spi_control_port_irq_from_sa),
      .sys_clk_freq_s1_irq_from_sa                                                         (sys_clk_freq_s1_irq_from_sa),
      .uart_0_s1_irq_from_sa                                                               (uart_0_s1_irq_from_sa)
    );

  cpu_linux_instruction_master_arbitrator the_cpu_linux_instruction_master
    (
      .Medipix_sopc_burst_0_upstream_readdata_from_sa                                            (Medipix_sopc_burst_0_upstream_readdata_from_sa),
      .Medipix_sopc_burst_0_upstream_waitrequest_from_sa                                         (Medipix_sopc_burst_0_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_4_upstream_readdata_from_sa                                            (Medipix_sopc_burst_4_upstream_readdata_from_sa),
      .Medipix_sopc_burst_4_upstream_waitrequest_from_sa                                         (Medipix_sopc_burst_4_upstream_waitrequest_from_sa),
      .Medipix_sopc_burst_6_upstream_readdata_from_sa                                            (Medipix_sopc_burst_6_upstream_readdata_from_sa),
      .Medipix_sopc_burst_6_upstream_waitrequest_from_sa                                         (Medipix_sopc_burst_6_upstream_waitrequest_from_sa),
      .clk                                                                                       (ram_aux_half_rate_clk_out),
      .cpu_linux_instruction_master_address                                                      (cpu_linux_instruction_master_address),
      .cpu_linux_instruction_master_address_to_slave                                             (cpu_linux_instruction_master_address_to_slave),
      .cpu_linux_instruction_master_burstcount                                                   (cpu_linux_instruction_master_burstcount),
      .cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream                        (cpu_linux_instruction_master_granted_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream                        (cpu_linux_instruction_master_granted_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream                        (cpu_linux_instruction_master_granted_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_latency_counter                                              (cpu_linux_instruction_master_latency_counter),
      .cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream              (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream              (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream              (cpu_linux_instruction_master_qualified_request_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_read                                                         (cpu_linux_instruction_master_read),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream                (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_0_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream                (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_4_upstream_shift_register),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream                (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register (cpu_linux_instruction_master_read_data_valid_Medipix_sopc_burst_6_upstream_shift_register),
      .cpu_linux_instruction_master_readdata                                                     (cpu_linux_instruction_master_readdata),
      .cpu_linux_instruction_master_readdatavalid                                                (cpu_linux_instruction_master_readdatavalid),
      .cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream                       (cpu_linux_instruction_master_requests_Medipix_sopc_burst_0_upstream),
      .cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream                       (cpu_linux_instruction_master_requests_Medipix_sopc_burst_4_upstream),
      .cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream                       (cpu_linux_instruction_master_requests_Medipix_sopc_burst_6_upstream),
      .cpu_linux_instruction_master_waitrequest                                                  (cpu_linux_instruction_master_waitrequest),
      .d1_Medipix_sopc_burst_0_upstream_end_xfer                                                 (d1_Medipix_sopc_burst_0_upstream_end_xfer),
      .d1_Medipix_sopc_burst_4_upstream_end_xfer                                                 (d1_Medipix_sopc_burst_4_upstream_end_xfer),
      .d1_Medipix_sopc_burst_6_upstream_end_xfer                                                 (d1_Medipix_sopc_burst_6_upstream_end_xfer),
      .reset_n                                                                                   (ram_aux_half_rate_clk_out_reset_n)
    );

  cpu_linux the_cpu_linux
    (
      .clk                                   (ram_aux_half_rate_clk_out),
      .d_address                             (cpu_linux_data_master_address),
      .d_burstcount                          (cpu_linux_data_master_burstcount),
      .d_byteenable                          (cpu_linux_data_master_byteenable),
      .d_irq                                 (cpu_linux_data_master_irq),
      .d_read                                (cpu_linux_data_master_read),
      .d_readdata                            (cpu_linux_data_master_readdata),
      .d_readdatavalid                       (cpu_linux_data_master_readdatavalid),
      .d_waitrequest                         (cpu_linux_data_master_waitrequest),
      .d_write                               (cpu_linux_data_master_write),
      .d_writedata                           (cpu_linux_data_master_writedata),
      .i_address                             (cpu_linux_instruction_master_address),
      .i_burstcount                          (cpu_linux_instruction_master_burstcount),
      .i_read                                (cpu_linux_instruction_master_read),
      .i_readdata                            (cpu_linux_instruction_master_readdata),
      .i_readdatavalid                       (cpu_linux_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_linux_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_linux_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_linux_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_linux_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_linux_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_linux_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_linux_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_linux_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_linux_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_linux_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_linux_jtag_debug_module_writedata),
      .reset_n                               (cpu_linux_jtag_debug_module_reset_n)
    );

  epcs_controller_epcs_control_port_arbitrator the_epcs_controller_epcs_control_port
    (
      .Medipix_sopc_burst_6_downstream_address_to_slave                                    (Medipix_sopc_burst_6_downstream_address_to_slave),
      .Medipix_sopc_burst_6_downstream_arbitrationshare                                    (Medipix_sopc_burst_6_downstream_arbitrationshare),
      .Medipix_sopc_burst_6_downstream_burstcount                                          (Medipix_sopc_burst_6_downstream_burstcount),
      .Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port           (Medipix_sopc_burst_6_downstream_granted_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_latency_counter                                     (Medipix_sopc_burst_6_downstream_latency_counter),
      .Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port (Medipix_sopc_burst_6_downstream_qualified_request_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_read                                                (Medipix_sopc_burst_6_downstream_read),
      .Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port   (Medipix_sopc_burst_6_downstream_read_data_valid_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port          (Medipix_sopc_burst_6_downstream_requests_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_6_downstream_write                                               (Medipix_sopc_burst_6_downstream_write),
      .Medipix_sopc_burst_6_downstream_writedata                                           (Medipix_sopc_burst_6_downstream_writedata),
      .Medipix_sopc_burst_7_downstream_address_to_slave                                    (Medipix_sopc_burst_7_downstream_address_to_slave),
      .Medipix_sopc_burst_7_downstream_arbitrationshare                                    (Medipix_sopc_burst_7_downstream_arbitrationshare),
      .Medipix_sopc_burst_7_downstream_burstcount                                          (Medipix_sopc_burst_7_downstream_burstcount),
      .Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port           (Medipix_sopc_burst_7_downstream_granted_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_latency_counter                                     (Medipix_sopc_burst_7_downstream_latency_counter),
      .Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port (Medipix_sopc_burst_7_downstream_qualified_request_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_read                                                (Medipix_sopc_burst_7_downstream_read),
      .Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port   (Medipix_sopc_burst_7_downstream_read_data_valid_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port          (Medipix_sopc_burst_7_downstream_requests_epcs_controller_epcs_control_port),
      .Medipix_sopc_burst_7_downstream_write                                               (Medipix_sopc_burst_7_downstream_write),
      .Medipix_sopc_burst_7_downstream_writedata                                           (Medipix_sopc_burst_7_downstream_writedata),
      .clk                                                                                 (ram_aux_half_rate_clk_out),
      .d1_epcs_controller_epcs_control_port_end_xfer                                       (d1_epcs_controller_epcs_control_port_end_xfer),
      .epcs_controller_epcs_control_port_address                                           (epcs_controller_epcs_control_port_address),
      .epcs_controller_epcs_control_port_chipselect                                        (epcs_controller_epcs_control_port_chipselect),
      .epcs_controller_epcs_control_port_dataavailable                                     (epcs_controller_epcs_control_port_dataavailable),
      .epcs_controller_epcs_control_port_dataavailable_from_sa                             (epcs_controller_epcs_control_port_dataavailable_from_sa),
      .epcs_controller_epcs_control_port_endofpacket                                       (epcs_controller_epcs_control_port_endofpacket),
      .epcs_controller_epcs_control_port_endofpacket_from_sa                               (epcs_controller_epcs_control_port_endofpacket_from_sa),
      .epcs_controller_epcs_control_port_irq                                               (epcs_controller_epcs_control_port_irq),
      .epcs_controller_epcs_control_port_irq_from_sa                                       (epcs_controller_epcs_control_port_irq_from_sa),
      .epcs_controller_epcs_control_port_read_n                                            (epcs_controller_epcs_control_port_read_n),
      .epcs_controller_epcs_control_port_readdata                                          (epcs_controller_epcs_control_port_readdata),
      .epcs_controller_epcs_control_port_readdata_from_sa                                  (epcs_controller_epcs_control_port_readdata_from_sa),
      .epcs_controller_epcs_control_port_readyfordata                                      (epcs_controller_epcs_control_port_readyfordata),
      .epcs_controller_epcs_control_port_readyfordata_from_sa                              (epcs_controller_epcs_control_port_readyfordata_from_sa),
      .epcs_controller_epcs_control_port_reset_n                                           (epcs_controller_epcs_control_port_reset_n),
      .epcs_controller_epcs_control_port_write_n                                           (epcs_controller_epcs_control_port_write_n),
      .epcs_controller_epcs_control_port_writedata                                         (epcs_controller_epcs_control_port_writedata),
      .reset_n                                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  epcs_controller the_epcs_controller
    (
      .address       (epcs_controller_epcs_control_port_address),
      .chipselect    (epcs_controller_epcs_control_port_chipselect),
      .clk           (ram_aux_half_rate_clk_out),
      .data0         (data0_to_the_epcs_controller),
      .dataavailable (epcs_controller_epcs_control_port_dataavailable),
      .dclk          (dclk_from_the_epcs_controller),
      .endofpacket   (epcs_controller_epcs_control_port_endofpacket),
      .irq           (epcs_controller_epcs_control_port_irq),
      .read_n        (epcs_controller_epcs_control_port_read_n),
      .readdata      (epcs_controller_epcs_control_port_readdata),
      .readyfordata  (epcs_controller_epcs_control_port_readyfordata),
      .reset_n       (epcs_controller_epcs_control_port_reset_n),
      .sce           (sce_from_the_epcs_controller),
      .sdo           (sdo_from_the_epcs_controller),
      .write_n       (epcs_controller_epcs_control_port_write_n),
      .writedata     (epcs_controller_epcs_control_port_writedata)
    );

  igor_mac_control_port_arbitrator the_igor_mac_control_port
    (
      .Medipix_sopc_burst_8_downstream_address_to_slave                        (Medipix_sopc_burst_8_downstream_address_to_slave),
      .Medipix_sopc_burst_8_downstream_arbitrationshare                        (Medipix_sopc_burst_8_downstream_arbitrationshare),
      .Medipix_sopc_burst_8_downstream_burstcount                              (Medipix_sopc_burst_8_downstream_burstcount),
      .Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port           (Medipix_sopc_burst_8_downstream_granted_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_latency_counter                         (Medipix_sopc_burst_8_downstream_latency_counter),
      .Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port (Medipix_sopc_burst_8_downstream_qualified_request_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_read                                    (Medipix_sopc_burst_8_downstream_read),
      .Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port   (Medipix_sopc_burst_8_downstream_read_data_valid_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port          (Medipix_sopc_burst_8_downstream_requests_igor_mac_control_port),
      .Medipix_sopc_burst_8_downstream_write                                   (Medipix_sopc_burst_8_downstream_write),
      .Medipix_sopc_burst_8_downstream_writedata                               (Medipix_sopc_burst_8_downstream_writedata),
      .clk                                                                     (ram_aux_half_rate_clk_out),
      .d1_igor_mac_control_port_end_xfer                                       (d1_igor_mac_control_port_end_xfer),
      .igor_mac_control_port_address                                           (igor_mac_control_port_address),
      .igor_mac_control_port_chipselect                                        (igor_mac_control_port_chipselect),
      .igor_mac_control_port_irq                                               (igor_mac_control_port_irq),
      .igor_mac_control_port_irq_from_sa                                       (igor_mac_control_port_irq_from_sa),
      .igor_mac_control_port_read                                              (igor_mac_control_port_read),
      .igor_mac_control_port_readdata                                          (igor_mac_control_port_readdata),
      .igor_mac_control_port_readdata_from_sa                                  (igor_mac_control_port_readdata_from_sa),
      .igor_mac_control_port_reset                                             (igor_mac_control_port_reset),
      .igor_mac_control_port_waitrequest_n                                     (igor_mac_control_port_waitrequest_n),
      .igor_mac_control_port_waitrequest_n_from_sa                             (igor_mac_control_port_waitrequest_n_from_sa),
      .igor_mac_control_port_write                                             (igor_mac_control_port_write),
      .igor_mac_control_port_writedata                                         (igor_mac_control_port_writedata),
      .reset_n                                                                 (ram_aux_half_rate_clk_out_reset_n)
    );

  igor_mac_rx_master_arbitrator the_igor_mac_rx_master
    (
      .clk                                                    (ram_aux_half_rate_clk_out),
      .clock_crossing_s1_waitrequest_from_sa                  (clock_crossing_s1_waitrequest_from_sa),
      .d1_clock_crossing_s1_end_xfer                          (d1_clock_crossing_s1_end_xfer),
      .igor_mac_rx_master_address                             (igor_mac_rx_master_address),
      .igor_mac_rx_master_address_to_slave                    (igor_mac_rx_master_address_to_slave),
      .igor_mac_rx_master_byteenable                          (igor_mac_rx_master_byteenable),
      .igor_mac_rx_master_granted_clock_crossing_s1           (igor_mac_rx_master_granted_clock_crossing_s1),
      .igor_mac_rx_master_qualified_request_clock_crossing_s1 (igor_mac_rx_master_qualified_request_clock_crossing_s1),
      .igor_mac_rx_master_requests_clock_crossing_s1          (igor_mac_rx_master_requests_clock_crossing_s1),
      .igor_mac_rx_master_waitrequest                         (igor_mac_rx_master_waitrequest),
      .igor_mac_rx_master_write                               (igor_mac_rx_master_write),
      .igor_mac_rx_master_writedata                           (igor_mac_rx_master_writedata),
      .reset_n                                                (ram_aux_half_rate_clk_out_reset_n)
    );

  igor_mac_tx_master_arbitrator the_igor_mac_tx_master
    (
      .clk                                                                 (ram_aux_half_rate_clk_out),
      .clock_crossing_s1_readdata_from_sa                                  (clock_crossing_s1_readdata_from_sa),
      .clock_crossing_s1_waitrequest_from_sa                               (clock_crossing_s1_waitrequest_from_sa),
      .d1_clock_crossing_s1_end_xfer                                       (d1_clock_crossing_s1_end_xfer),
      .igor_mac_tx_master_address                                          (igor_mac_tx_master_address),
      .igor_mac_tx_master_address_to_slave                                 (igor_mac_tx_master_address_to_slave),
      .igor_mac_tx_master_granted_clock_crossing_s1                        (igor_mac_tx_master_granted_clock_crossing_s1),
      .igor_mac_tx_master_latency_counter                                  (igor_mac_tx_master_latency_counter),
      .igor_mac_tx_master_qualified_request_clock_crossing_s1              (igor_mac_tx_master_qualified_request_clock_crossing_s1),
      .igor_mac_tx_master_read                                             (igor_mac_tx_master_read),
      .igor_mac_tx_master_read_data_valid_clock_crossing_s1                (igor_mac_tx_master_read_data_valid_clock_crossing_s1),
      .igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register (igor_mac_tx_master_read_data_valid_clock_crossing_s1_shift_register),
      .igor_mac_tx_master_readdata                                         (igor_mac_tx_master_readdata),
      .igor_mac_tx_master_readdatavalid                                    (igor_mac_tx_master_readdatavalid),
      .igor_mac_tx_master_requests_clock_crossing_s1                       (igor_mac_tx_master_requests_clock_crossing_s1),
      .igor_mac_tx_master_waitrequest                                      (igor_mac_tx_master_waitrequest),
      .reset_n                                                             (ram_aux_half_rate_clk_out_reset_n)
    );

  igor_mac the_igor_mac
    (
      .av_address          (igor_mac_control_port_address),
      .av_chipselect       (igor_mac_control_port_chipselect),
      .av_clk              (ram_aux_half_rate_clk_out),
      .av_irq              (igor_mac_control_port_irq),
      .av_read             (igor_mac_control_port_read),
      .av_readdata         (igor_mac_control_port_readdata),
      .av_reset            (igor_mac_control_port_reset),
      .av_rx_address       (igor_mac_rx_master_address),
      .av_rx_byteenable    (igor_mac_rx_master_byteenable),
      .av_rx_waitrequest   (igor_mac_rx_master_waitrequest),
      .av_rx_write         (igor_mac_rx_master_write),
      .av_rx_writedata     (igor_mac_rx_master_writedata),
      .av_tx_address       (igor_mac_tx_master_address),
      .av_tx_read          (igor_mac_tx_master_read),
      .av_tx_readdata      (igor_mac_tx_master_readdata),
      .av_tx_readdatavalid (igor_mac_tx_master_readdatavalid),
      .av_tx_waitrequest   (igor_mac_tx_master_waitrequest),
      .av_waitrequest_n    (igor_mac_control_port_waitrequest_n),
      .av_write            (igor_mac_control_port_write),
      .av_writedata        (igor_mac_control_port_writedata),
      .mcoll_pad_i         (mcoll_pad_i_to_the_igor_mac),
      .mcrs_pad_i          (mcrs_pad_i_to_the_igor_mac),
      .md_pad_i            (md_pad_i_to_the_igor_mac),
      .md_pad_o            (md_pad_o_from_the_igor_mac),
      .md_padoe_o          (md_padoe_o_from_the_igor_mac),
      .mdc_pad_o           (mdc_pad_o_from_the_igor_mac),
      .mrx_clk_pad_i       (mrx_clk_pad_i_to_the_igor_mac),
      .mrxd_pad_i          (mrxd_pad_i_to_the_igor_mac),
      .mrxdv_pad_i         (mrxdv_pad_i_to_the_igor_mac),
      .mrxerr_pad_i        (mrxerr_pad_i_to_the_igor_mac),
      .mtx_clk_pad_i       (mtx_clk_pad_i_to_the_igor_mac),
      .mtxd_pad_o          (mtxd_pad_o_from_the_igor_mac),
      .mtxen_pad_o         (mtxen_pad_o_from_the_igor_mac),
      .mtxerr_pad_o        (mtxerr_pad_o_from_the_igor_mac)
    );

  jtag_uart_0_avalon_jtag_slave_arbitrator the_jtag_uart_0_avalon_jtag_slave
    (
      .Medipix_sopc_burst_2_downstream_address_to_slave                                (Medipix_sopc_burst_2_downstream_address_to_slave),
      .Medipix_sopc_burst_2_downstream_arbitrationshare                                (Medipix_sopc_burst_2_downstream_arbitrationshare),
      .Medipix_sopc_burst_2_downstream_burstcount                                      (Medipix_sopc_burst_2_downstream_burstcount),
      .Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave           (Medipix_sopc_burst_2_downstream_granted_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_latency_counter                                 (Medipix_sopc_burst_2_downstream_latency_counter),
      .Medipix_sopc_burst_2_downstream_nativeaddress                                   (Medipix_sopc_burst_2_downstream_nativeaddress),
      .Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave (Medipix_sopc_burst_2_downstream_qualified_request_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_read                                            (Medipix_sopc_burst_2_downstream_read),
      .Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave   (Medipix_sopc_burst_2_downstream_read_data_valid_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave          (Medipix_sopc_burst_2_downstream_requests_jtag_uart_0_avalon_jtag_slave),
      .Medipix_sopc_burst_2_downstream_write                                           (Medipix_sopc_burst_2_downstream_write),
      .Medipix_sopc_burst_2_downstream_writedata                                       (Medipix_sopc_burst_2_downstream_writedata),
      .clk                                                                             (ram_aux_half_rate_clk_out),
      .d1_jtag_uart_0_avalon_jtag_slave_end_xfer                                       (d1_jtag_uart_0_avalon_jtag_slave_end_xfer),
      .jtag_uart_0_avalon_jtag_slave_address                                           (jtag_uart_0_avalon_jtag_slave_address),
      .jtag_uart_0_avalon_jtag_slave_chipselect                                        (jtag_uart_0_avalon_jtag_slave_chipselect),
      .jtag_uart_0_avalon_jtag_slave_dataavailable                                     (jtag_uart_0_avalon_jtag_slave_dataavailable),
      .jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa                             (jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_0_avalon_jtag_slave_irq                                               (jtag_uart_0_avalon_jtag_slave_irq),
      .jtag_uart_0_avalon_jtag_slave_irq_from_sa                                       (jtag_uart_0_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_0_avalon_jtag_slave_read_n                                            (jtag_uart_0_avalon_jtag_slave_read_n),
      .jtag_uart_0_avalon_jtag_slave_readdata                                          (jtag_uart_0_avalon_jtag_slave_readdata),
      .jtag_uart_0_avalon_jtag_slave_readdata_from_sa                                  (jtag_uart_0_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_readyfordata                                      (jtag_uart_0_avalon_jtag_slave_readyfordata),
      .jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa                              (jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_reset_n                                           (jtag_uart_0_avalon_jtag_slave_reset_n),
      .jtag_uart_0_avalon_jtag_slave_waitrequest                                       (jtag_uart_0_avalon_jtag_slave_waitrequest),
      .jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa                               (jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_0_avalon_jtag_slave_write_n                                           (jtag_uart_0_avalon_jtag_slave_write_n),
      .jtag_uart_0_avalon_jtag_slave_writedata                                         (jtag_uart_0_avalon_jtag_slave_writedata),
      .reset_n                                                                         (ram_aux_half_rate_clk_out_reset_n)
    );

  jtag_uart_0 the_jtag_uart_0
    (
      .av_address     (jtag_uart_0_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_0_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_0_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_0_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_0_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_0_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_0_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_0_avalon_jtag_slave_writedata),
      .clk            (ram_aux_half_rate_clk_out),
      .dataavailable  (jtag_uart_0_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_0_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_0_avalon_jtag_slave_reset_n)
    );

  ram_s1_arbitrator the_ram_s1
    (
      .clk                                                     (ram_phy_clk_out),
      .clock_crossing_m1_address_to_slave                      (clock_crossing_m1_address_to_slave),
      .clock_crossing_m1_byteenable                            (clock_crossing_m1_byteenable),
      .clock_crossing_m1_granted_ram_s1                        (clock_crossing_m1_granted_ram_s1),
      .clock_crossing_m1_latency_counter                       (clock_crossing_m1_latency_counter),
      .clock_crossing_m1_qualified_request_ram_s1              (clock_crossing_m1_qualified_request_ram_s1),
      .clock_crossing_m1_read                                  (clock_crossing_m1_read),
      .clock_crossing_m1_read_data_valid_ram_s1                (clock_crossing_m1_read_data_valid_ram_s1),
      .clock_crossing_m1_read_data_valid_ram_s1_shift_register (clock_crossing_m1_read_data_valid_ram_s1_shift_register),
      .clock_crossing_m1_requests_ram_s1                       (clock_crossing_m1_requests_ram_s1),
      .clock_crossing_m1_write                                 (clock_crossing_m1_write),
      .clock_crossing_m1_writedata                             (clock_crossing_m1_writedata),
      .d1_ram_s1_end_xfer                                      (d1_ram_s1_end_xfer),
      .ram_s1_address                                          (ram_s1_address),
      .ram_s1_beginbursttransfer                               (ram_s1_beginbursttransfer),
      .ram_s1_burstcount                                       (ram_s1_burstcount),
      .ram_s1_byteenable                                       (ram_s1_byteenable),
      .ram_s1_read                                             (ram_s1_read),
      .ram_s1_readdata                                         (ram_s1_readdata),
      .ram_s1_readdata_from_sa                                 (ram_s1_readdata_from_sa),
      .ram_s1_readdatavalid                                    (ram_s1_readdatavalid),
      .ram_s1_resetrequest_n                                   (ram_s1_resetrequest_n),
      .ram_s1_resetrequest_n_from_sa                           (ram_s1_resetrequest_n_from_sa),
      .ram_s1_waitrequest_n                                    (ram_s1_waitrequest_n),
      .ram_s1_waitrequest_n_from_sa                            (ram_s1_waitrequest_n_from_sa),
      .ram_s1_write                                            (ram_s1_write),
      .ram_s1_writedata                                        (ram_s1_writedata),
      .reset_n                                                 (ram_phy_clk_out_reset_n)
    );

  //ram_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  assign ram_aux_full_rate_clk_out = out_clk_ram_aux_full_rate_clk;

  //ram_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  assign ram_aux_half_rate_clk_out = out_clk_ram_aux_half_rate_clk;

  //ram_phy_clk_out out_clk assignment, which is an e_assign
  assign ram_phy_clk_out = out_clk_ram_phy_clk;

  //reset is asserted asynchronously and deasserted synchronously
  Medipix_sopc_reset_clk_125_domain_synch_module Medipix_sopc_reset_clk_125_domain_synch
    (
      .clk      (clk_125),
      .data_in  (1'b1),
      .data_out (clk_125_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    0 |
    cpu_linux_jtag_debug_module_resetrequest_from_sa |
    cpu_linux_jtag_debug_module_resetrequest_from_sa |
    0 |
    ~ram_s1_resetrequest_n_from_sa |
    ~ram_s1_resetrequest_n_from_sa);

  ram the_ram
    (
      .aux_full_rate_clk (out_clk_ram_aux_full_rate_clk),
      .aux_half_rate_clk (out_clk_ram_aux_half_rate_clk),
      .global_reset_n    (global_reset_n_to_the_ram),
      .local_address     (ram_s1_address),
      .local_be          (ram_s1_byteenable),
      .local_burstbegin  (ram_s1_beginbursttransfer),
      .local_init_done   (local_init_done_from_the_ram),
      .local_rdata       (ram_s1_readdata),
      .local_rdata_valid (ram_s1_readdatavalid),
      .local_read_req    (ram_s1_read),
      .local_ready       (ram_s1_waitrequest_n),
      .local_refresh_ack (local_refresh_ack_from_the_ram),
      .local_size        (ram_s1_burstcount),
      .local_wdata       (ram_s1_writedata),
      .local_wdata_req   (local_wdata_req_from_the_ram),
      .local_write_req   (ram_s1_write),
      .mem_addr          (mem_addr_from_the_ram),
      .mem_ba            (mem_ba_from_the_ram),
      .mem_cas_n         (mem_cas_n_from_the_ram),
      .mem_cke           (mem_cke_from_the_ram),
      .mem_clk           (mem_clk_to_and_from_the_ram),
      .mem_clk_n         (mem_clk_n_to_and_from_the_ram),
      .mem_cs_n          (mem_cs_n_from_the_ram),
      .mem_dm            (mem_dm_from_the_ram),
      .mem_dq            (mem_dq_to_and_from_the_ram),
      .mem_dqs           (mem_dqs_to_and_from_the_ram),
      .mem_odt           (mem_odt_from_the_ram),
      .mem_ras_n         (mem_ras_n_from_the_ram),
      .mem_we_n          (mem_we_n_from_the_ram),
      .phy_clk           (out_clk_ram_phy_clk),
      .pll_ref_clk       (clk_125),
      .reset_phy_clk_n   (reset_phy_clk_n_from_the_ram),
      .reset_request_n   (ram_s1_resetrequest_n),
      .soft_reset_n      (clk_125_reset_n)
    );

  spi_0_spi_control_port_arbitrator the_spi_0_spi_control_port
    (
      .Medipix_sopc_burst_10_downstream_address_to_slave                         (Medipix_sopc_burst_10_downstream_address_to_slave),
      .Medipix_sopc_burst_10_downstream_arbitrationshare                         (Medipix_sopc_burst_10_downstream_arbitrationshare),
      .Medipix_sopc_burst_10_downstream_burstcount                               (Medipix_sopc_burst_10_downstream_burstcount),
      .Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port           (Medipix_sopc_burst_10_downstream_granted_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_latency_counter                          (Medipix_sopc_burst_10_downstream_latency_counter),
      .Medipix_sopc_burst_10_downstream_nativeaddress                            (Medipix_sopc_burst_10_downstream_nativeaddress),
      .Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port (Medipix_sopc_burst_10_downstream_qualified_request_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_read                                     (Medipix_sopc_burst_10_downstream_read),
      .Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port   (Medipix_sopc_burst_10_downstream_read_data_valid_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port          (Medipix_sopc_burst_10_downstream_requests_spi_0_spi_control_port),
      .Medipix_sopc_burst_10_downstream_write                                    (Medipix_sopc_burst_10_downstream_write),
      .Medipix_sopc_burst_10_downstream_writedata                                (Medipix_sopc_burst_10_downstream_writedata),
      .clk                                                                       (ram_aux_half_rate_clk_out),
      .d1_spi_0_spi_control_port_end_xfer                                        (d1_spi_0_spi_control_port_end_xfer),
      .reset_n                                                                   (ram_aux_half_rate_clk_out_reset_n),
      .spi_0_spi_control_port_address                                            (spi_0_spi_control_port_address),
      .spi_0_spi_control_port_chipselect                                         (spi_0_spi_control_port_chipselect),
      .spi_0_spi_control_port_dataavailable                                      (spi_0_spi_control_port_dataavailable),
      .spi_0_spi_control_port_dataavailable_from_sa                              (spi_0_spi_control_port_dataavailable_from_sa),
      .spi_0_spi_control_port_endofpacket                                        (spi_0_spi_control_port_endofpacket),
      .spi_0_spi_control_port_endofpacket_from_sa                                (spi_0_spi_control_port_endofpacket_from_sa),
      .spi_0_spi_control_port_irq                                                (spi_0_spi_control_port_irq),
      .spi_0_spi_control_port_irq_from_sa                                        (spi_0_spi_control_port_irq_from_sa),
      .spi_0_spi_control_port_read_n                                             (spi_0_spi_control_port_read_n),
      .spi_0_spi_control_port_readdata                                           (spi_0_spi_control_port_readdata),
      .spi_0_spi_control_port_readdata_from_sa                                   (spi_0_spi_control_port_readdata_from_sa),
      .spi_0_spi_control_port_readyfordata                                       (spi_0_spi_control_port_readyfordata),
      .spi_0_spi_control_port_readyfordata_from_sa                               (spi_0_spi_control_port_readyfordata_from_sa),
      .spi_0_spi_control_port_reset_n                                            (spi_0_spi_control_port_reset_n),
      .spi_0_spi_control_port_write_n                                            (spi_0_spi_control_port_write_n),
      .spi_0_spi_control_port_writedata                                          (spi_0_spi_control_port_writedata)
    );

  spi_0 the_spi_0
    (
      .MISO          (MISO_to_the_spi_0),
      .MOSI          (MOSI_from_the_spi_0),
      .SCLK          (SCLK_from_the_spi_0),
      .SS_n          (SS_n_from_the_spi_0),
      .clk           (ram_aux_half_rate_clk_out),
      .data_from_cpu (spi_0_spi_control_port_writedata),
      .data_to_cpu   (spi_0_spi_control_port_readdata),
      .dataavailable (spi_0_spi_control_port_dataavailable),
      .endofpacket   (spi_0_spi_control_port_endofpacket),
      .irq           (spi_0_spi_control_port_irq),
      .mem_addr      (spi_0_spi_control_port_address),
      .read_n        (spi_0_spi_control_port_read_n),
      .readyfordata  (spi_0_spi_control_port_readyfordata),
      .reset_n       (spi_0_spi_control_port_reset_n),
      .spi_select    (spi_0_spi_control_port_chipselect),
      .write_n       (spi_0_spi_control_port_write_n)
    );

  sys_clk_freq_s1_arbitrator the_sys_clk_freq_s1
    (
      .Medipix_sopc_burst_3_downstream_address_to_slave                  (Medipix_sopc_burst_3_downstream_address_to_slave),
      .Medipix_sopc_burst_3_downstream_arbitrationshare                  (Medipix_sopc_burst_3_downstream_arbitrationshare),
      .Medipix_sopc_burst_3_downstream_burstcount                        (Medipix_sopc_burst_3_downstream_burstcount),
      .Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1           (Medipix_sopc_burst_3_downstream_granted_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_latency_counter                   (Medipix_sopc_burst_3_downstream_latency_counter),
      .Medipix_sopc_burst_3_downstream_nativeaddress                     (Medipix_sopc_burst_3_downstream_nativeaddress),
      .Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1 (Medipix_sopc_burst_3_downstream_qualified_request_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_read                              (Medipix_sopc_burst_3_downstream_read),
      .Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1   (Medipix_sopc_burst_3_downstream_read_data_valid_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1          (Medipix_sopc_burst_3_downstream_requests_sys_clk_freq_s1),
      .Medipix_sopc_burst_3_downstream_write                             (Medipix_sopc_burst_3_downstream_write),
      .Medipix_sopc_burst_3_downstream_writedata                         (Medipix_sopc_burst_3_downstream_writedata),
      .clk                                                               (ram_aux_half_rate_clk_out),
      .d1_sys_clk_freq_s1_end_xfer                                       (d1_sys_clk_freq_s1_end_xfer),
      .reset_n                                                           (ram_aux_half_rate_clk_out_reset_n),
      .sys_clk_freq_s1_address                                           (sys_clk_freq_s1_address),
      .sys_clk_freq_s1_chipselect                                        (sys_clk_freq_s1_chipselect),
      .sys_clk_freq_s1_irq                                               (sys_clk_freq_s1_irq),
      .sys_clk_freq_s1_irq_from_sa                                       (sys_clk_freq_s1_irq_from_sa),
      .sys_clk_freq_s1_readdata                                          (sys_clk_freq_s1_readdata),
      .sys_clk_freq_s1_readdata_from_sa                                  (sys_clk_freq_s1_readdata_from_sa),
      .sys_clk_freq_s1_reset_n                                           (sys_clk_freq_s1_reset_n),
      .sys_clk_freq_s1_write_n                                           (sys_clk_freq_s1_write_n),
      .sys_clk_freq_s1_writedata                                         (sys_clk_freq_s1_writedata)
    );

  sys_clk_freq the_sys_clk_freq
    (
      .address    (sys_clk_freq_s1_address),
      .chipselect (sys_clk_freq_s1_chipselect),
      .clk        (ram_aux_half_rate_clk_out),
      .irq        (sys_clk_freq_s1_irq),
      .readdata   (sys_clk_freq_s1_readdata),
      .reset_n    (sys_clk_freq_s1_reset_n),
      .write_n    (sys_clk_freq_s1_write_n),
      .writedata  (sys_clk_freq_s1_writedata)
    );

  tx_table_avalon_slave_0_arbitrator the_tx_table_avalon_slave_0
    (
      .Medipix_sopc_burst_9_downstream_address_to_slave                          (Medipix_sopc_burst_9_downstream_address_to_slave),
      .Medipix_sopc_burst_9_downstream_arbitrationshare                          (Medipix_sopc_burst_9_downstream_arbitrationshare),
      .Medipix_sopc_burst_9_downstream_burstcount                                (Medipix_sopc_burst_9_downstream_burstcount),
      .Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0           (Medipix_sopc_burst_9_downstream_granted_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_latency_counter                           (Medipix_sopc_burst_9_downstream_latency_counter),
      .Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0 (Medipix_sopc_burst_9_downstream_qualified_request_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_read                                      (Medipix_sopc_burst_9_downstream_read),
      .Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0   (Medipix_sopc_burst_9_downstream_read_data_valid_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0          (Medipix_sopc_burst_9_downstream_requests_tx_table_avalon_slave_0),
      .Medipix_sopc_burst_9_downstream_write                                     (Medipix_sopc_burst_9_downstream_write),
      .Medipix_sopc_burst_9_downstream_writedata                                 (Medipix_sopc_burst_9_downstream_writedata),
      .clk                                                                       (ram_aux_half_rate_clk_out),
      .d1_tx_table_avalon_slave_0_end_xfer                                       (d1_tx_table_avalon_slave_0_end_xfer),
      .reset_n                                                                   (ram_aux_half_rate_clk_out_reset_n),
      .tx_table_avalon_slave_0_address                                           (tx_table_avalon_slave_0_address),
      .tx_table_avalon_slave_0_chipselect                                        (tx_table_avalon_slave_0_chipselect),
      .tx_table_avalon_slave_0_read                                              (tx_table_avalon_slave_0_read),
      .tx_table_avalon_slave_0_readdata                                          (tx_table_avalon_slave_0_readdata),
      .tx_table_avalon_slave_0_readdata_from_sa                                  (tx_table_avalon_slave_0_readdata_from_sa),
      .tx_table_avalon_slave_0_reset_n                                           (tx_table_avalon_slave_0_reset_n),
      .tx_table_avalon_slave_0_write                                             (tx_table_avalon_slave_0_write),
      .tx_table_avalon_slave_0_writedata                                         (tx_table_avalon_slave_0_writedata)
    );

  tx_table the_tx_table
    (
      .address    (tx_table_avalon_slave_0_address),
      .chipselect (tx_table_avalon_slave_0_chipselect),
      .clk        (ram_aux_half_rate_clk_out),
      .clock_vhdl (clock_vhdl_to_the_tx_table),
      .in_Nreset  (in_Nreset_to_the_tx_table),
      .info_out   (info_out_from_the_tx_table),
      .irq        (irq_from_the_tx_table),
      .out_data   (out_data_from_the_tx_table),
      .out_sync   (out_sync_from_the_tx_table),
      .out_valid  (out_valid_from_the_tx_table),
      .read       (tx_table_avalon_slave_0_read),
      .readdata   (tx_table_avalon_slave_0_readdata),
      .rst_n      (tx_table_avalon_slave_0_reset_n),
      .write      (tx_table_avalon_slave_0_write),
      .writedata  (tx_table_avalon_slave_0_writedata)
    );

  uart_0_s1_arbitrator the_uart_0_s1
    (
      .Medipix_sopc_burst_11_downstream_address_to_slave            (Medipix_sopc_burst_11_downstream_address_to_slave),
      .Medipix_sopc_burst_11_downstream_arbitrationshare            (Medipix_sopc_burst_11_downstream_arbitrationshare),
      .Medipix_sopc_burst_11_downstream_burstcount                  (Medipix_sopc_burst_11_downstream_burstcount),
      .Medipix_sopc_burst_11_downstream_granted_uart_0_s1           (Medipix_sopc_burst_11_downstream_granted_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_latency_counter             (Medipix_sopc_burst_11_downstream_latency_counter),
      .Medipix_sopc_burst_11_downstream_nativeaddress               (Medipix_sopc_burst_11_downstream_nativeaddress),
      .Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1 (Medipix_sopc_burst_11_downstream_qualified_request_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_read                        (Medipix_sopc_burst_11_downstream_read),
      .Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1   (Medipix_sopc_burst_11_downstream_read_data_valid_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_requests_uart_0_s1          (Medipix_sopc_burst_11_downstream_requests_uart_0_s1),
      .Medipix_sopc_burst_11_downstream_write                       (Medipix_sopc_burst_11_downstream_write),
      .Medipix_sopc_burst_11_downstream_writedata                   (Medipix_sopc_burst_11_downstream_writedata),
      .clk                                                          (ram_aux_half_rate_clk_out),
      .d1_uart_0_s1_end_xfer                                        (d1_uart_0_s1_end_xfer),
      .reset_n                                                      (ram_aux_half_rate_clk_out_reset_n),
      .uart_0_s1_address                                            (uart_0_s1_address),
      .uart_0_s1_begintransfer                                      (uart_0_s1_begintransfer),
      .uart_0_s1_chipselect                                         (uart_0_s1_chipselect),
      .uart_0_s1_dataavailable                                      (uart_0_s1_dataavailable),
      .uart_0_s1_dataavailable_from_sa                              (uart_0_s1_dataavailable_from_sa),
      .uart_0_s1_irq                                                (uart_0_s1_irq),
      .uart_0_s1_irq_from_sa                                        (uart_0_s1_irq_from_sa),
      .uart_0_s1_read_n                                             (uart_0_s1_read_n),
      .uart_0_s1_readdata                                           (uart_0_s1_readdata),
      .uart_0_s1_readdata_from_sa                                   (uart_0_s1_readdata_from_sa),
      .uart_0_s1_readyfordata                                       (uart_0_s1_readyfordata),
      .uart_0_s1_readyfordata_from_sa                               (uart_0_s1_readyfordata_from_sa),
      .uart_0_s1_reset_n                                            (uart_0_s1_reset_n),
      .uart_0_s1_write_n                                            (uart_0_s1_write_n),
      .uart_0_s1_writedata                                          (uart_0_s1_writedata)
    );

  uart_0 the_uart_0
    (
      .address       (uart_0_s1_address),
      .begintransfer (uart_0_s1_begintransfer),
      .chipselect    (uart_0_s1_chipselect),
      .clk           (ram_aux_half_rate_clk_out),
      .dataavailable (uart_0_s1_dataavailable),
      .irq           (uart_0_s1_irq),
      .read_n        (uart_0_s1_read_n),
      .readdata      (uart_0_s1_readdata),
      .readyfordata  (uart_0_s1_readyfordata),
      .reset_n       (uart_0_s1_reset_n),
      .rxd           (rxd_to_the_uart_0),
      .txd           (txd_from_the_uart_0),
      .write_n       (uart_0_s1_write_n),
      .writedata     (uart_0_s1_writedata)
    );

  //reset is asserted asynchronously and deasserted synchronously
  Medipix_sopc_reset_ram_aux_half_rate_clk_out_domain_synch_module Medipix_sopc_reset_ram_aux_half_rate_clk_out_domain_synch
    (
      .clk      (ram_aux_half_rate_clk_out),
      .data_in  (1'b1),
      .data_out (ram_aux_half_rate_clk_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  Medipix_sopc_reset_ram_phy_clk_out_domain_synch_module Medipix_sopc_reset_ram_phy_clk_out_domain_synch
    (
      .clk      (ram_phy_clk_out),
      .data_in  (1'b1),
      .data_out (ram_phy_clk_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //Medipix_sopc_burst_0_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign Medipix_sopc_burst_0_upstream_writedata = 0;

  //Medipix_sopc_burst_4_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign Medipix_sopc_burst_4_upstream_writedata = 0;

  //Medipix_sopc_burst_6_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign Medipix_sopc_burst_6_upstream_writedata = 0;

  //clock_crossing_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign clock_crossing_m1_endofpacket = 0;


endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "d:/altera/10.0/quartus/eda/sim_lib/altera_mf.v"
`include "d:/altera/10.0/quartus/eda/sim_lib/220model.v"
`include "d:/altera/10.0/quartus/eda/sim_lib/sgate.v"
`include "eth_ocm/eth_ocm.v"
`include "igor_mac.v"
// Modules/m_Txtable/txtable.vhd
// Modules/m_Txtable/avalon_wrdata.vhd
// Modules/m_Txtable/txdata_tovhdl.vhd
// Modules/m_Txtable/IP_ram_txtable.vhd
// tx_table.vhd
`include "Medipix_sopc_burst_0.v"
`include "clock_crossing.v"
`include "Medipix_sopc_burst_3.v"
`include "cpu_linux_test_bench.v"
`include "cpu_linux_mult_cell.v"
`include "cpu_linux_oci_test_bench.v"
`include "cpu_linux_jtag_debug_module_tck.v"
`include "cpu_linux_jtag_debug_module_sysclk.v"
`include "cpu_linux_jtag_debug_module_wrapper.v"
`include "cpu_linux.v"
`include "Medipix_sopc_burst_9.v"
`include "uart_0.v"
`include "Medipix_sopc_burst_4.v"
`include "spi_0.v"
`include "jtag_uart_0.v"
`include "sys_clk_freq.v"
`include "Medipix_sopc_burst_5.v"
`include "Medipix_sopc_burst_7.v"
`include "Medipix_sopc_burst_2.v"
`include "Medipix_sopc_burst_8.v"
`include "Medipix_sopc_burst_1.v"
`include "Medipix_sopc_burst_11.v"
`include "Medipix_sopc_burst_10.v"
`include "Medipix_sopc_burst_6.v"
`include "epcs_controller.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire             MISO_to_the_spi_0;
  wire             MOSI_from_the_spi_0;
  wire    [ 10: 0] Medipix_sopc_burst_0_downstream_nativeaddress;
  wire    [ 31: 0] Medipix_sopc_burst_0_upstream_writedata;
  wire             Medipix_sopc_burst_10_downstream_debugaccess;
  wire             Medipix_sopc_burst_11_downstream_debugaccess;
  wire    [ 10: 0] Medipix_sopc_burst_1_downstream_nativeaddress;
  wire             Medipix_sopc_burst_2_downstream_debugaccess;
  wire             Medipix_sopc_burst_3_downstream_debugaccess;
  wire             Medipix_sopc_burst_4_downstream_debugaccess;
  wire    [ 31: 0] Medipix_sopc_burst_4_upstream_writedata;
  wire             Medipix_sopc_burst_5_downstream_debugaccess;
  wire             Medipix_sopc_burst_6_downstream_debugaccess;
  wire    [ 10: 0] Medipix_sopc_burst_6_downstream_nativeaddress;
  wire    [ 31: 0] Medipix_sopc_burst_6_upstream_writedata;
  wire             Medipix_sopc_burst_7_downstream_debugaccess;
  wire    [ 10: 0] Medipix_sopc_burst_7_downstream_nativeaddress;
  wire             Medipix_sopc_burst_8_downstream_debugaccess;
  wire    [ 11: 0] Medipix_sopc_burst_8_downstream_nativeaddress;
  wire             Medipix_sopc_burst_9_downstream_debugaccess;
  wire    [  3: 0] Medipix_sopc_burst_9_downstream_nativeaddress;
  wire             SCLK_from_the_spi_0;
  wire    [  1: 0] SS_n_from_the_spi_0;
  wire             clk;
  reg              clk_125;
  wire             clock_crossing_m1_endofpacket;
  wire    [ 24: 0] clock_crossing_m1_nativeaddress;
  wire             clock_crossing_s1_endofpacket_from_sa;
  wire             clock_vhdl_to_the_tx_table;
  wire             data0_to_the_epcs_controller;
  wire             dclk_from_the_epcs_controller;
  wire             epcs_controller_epcs_control_port_dataavailable_from_sa;
  wire             epcs_controller_epcs_control_port_endofpacket_from_sa;
  wire             epcs_controller_epcs_control_port_readyfordata_from_sa;
  wire             global_reset_n_to_the_ram;
  wire             in_Nreset_to_the_tx_table;
  wire    [  7: 0] info_out_from_the_tx_table;
  wire             irq_from_the_tx_table;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  wire             local_init_done_from_the_ram;
  wire             local_refresh_ack_from_the_ram;
  wire             local_wdata_req_from_the_ram;
  wire             mcoll_pad_i_to_the_igor_mac;
  wire             mcrs_pad_i_to_the_igor_mac;
  wire             md_pad_i_to_the_igor_mac;
  wire             md_pad_o_from_the_igor_mac;
  wire             md_padoe_o_from_the_igor_mac;
  wire             mdc_pad_o_from_the_igor_mac;
  wire    [ 12: 0] mem_addr_from_the_ram;
  wire    [  2: 0] mem_ba_from_the_ram;
  wire             mem_cas_n_from_the_ram;
  wire             mem_cke_from_the_ram;
  wire             mem_clk_n_to_and_from_the_ram;
  wire             mem_clk_to_and_from_the_ram;
  wire             mem_cs_n_from_the_ram;
  wire    [  1: 0] mem_dm_from_the_ram;
  wire    [ 15: 0] mem_dq_to_and_from_the_ram;
  wire    [  1: 0] mem_dqs_to_and_from_the_ram;
  wire             mem_odt_from_the_ram;
  wire             mem_ras_n_from_the_ram;
  wire             mem_we_n_from_the_ram;
  wire             mrx_clk_pad_i_to_the_igor_mac;
  wire    [  3: 0] mrxd_pad_i_to_the_igor_mac;
  wire             mrxdv_pad_i_to_the_igor_mac;
  wire             mrxerr_pad_i_to_the_igor_mac;
  wire             mtx_clk_pad_i_to_the_igor_mac;
  wire    [  3: 0] mtxd_pad_o_from_the_igor_mac;
  wire             mtxen_pad_o_from_the_igor_mac;
  wire             mtxerr_pad_o_from_the_igor_mac;
  wire    [  7: 0] out_data_from_the_tx_table;
  wire             out_sync_from_the_tx_table;
  wire             out_valid_from_the_tx_table;
  wire             ram_aux_full_rate_clk_out;
  wire             ram_aux_half_rate_clk_out;
  wire             ram_phy_clk_out;
  reg              reset_n;
  wire             reset_phy_clk_n_from_the_ram;
  wire             rxd_to_the_uart_0;
  wire             sce_from_the_epcs_controller;
  wire             sdo_from_the_epcs_controller;
  wire             spi_0_spi_control_port_dataavailable_from_sa;
  wire             spi_0_spi_control_port_endofpacket_from_sa;
  wire             spi_0_spi_control_port_readyfordata_from_sa;
  wire             txd_from_the_uart_0;
  wire             uart_0_s1_dataavailable_from_sa;
  wire             uart_0_s1_readyfordata_from_sa;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  Medipix_sopc DUT
    (
      .MISO_to_the_spi_0              (MISO_to_the_spi_0),
      .MOSI_from_the_spi_0            (MOSI_from_the_spi_0),
      .SCLK_from_the_spi_0            (SCLK_from_the_spi_0),
      .SS_n_from_the_spi_0            (SS_n_from_the_spi_0),
      .clk_125                        (clk_125),
      .clock_vhdl_to_the_tx_table     (clock_vhdl_to_the_tx_table),
      .data0_to_the_epcs_controller   (data0_to_the_epcs_controller),
      .dclk_from_the_epcs_controller  (dclk_from_the_epcs_controller),
      .global_reset_n_to_the_ram      (global_reset_n_to_the_ram),
      .in_Nreset_to_the_tx_table      (in_Nreset_to_the_tx_table),
      .info_out_from_the_tx_table     (info_out_from_the_tx_table),
      .irq_from_the_tx_table          (irq_from_the_tx_table),
      .local_init_done_from_the_ram   (local_init_done_from_the_ram),
      .local_refresh_ack_from_the_ram (local_refresh_ack_from_the_ram),
      .local_wdata_req_from_the_ram   (local_wdata_req_from_the_ram),
      .mcoll_pad_i_to_the_igor_mac    (mcoll_pad_i_to_the_igor_mac),
      .mcrs_pad_i_to_the_igor_mac     (mcrs_pad_i_to_the_igor_mac),
      .md_pad_i_to_the_igor_mac       (md_pad_i_to_the_igor_mac),
      .md_pad_o_from_the_igor_mac     (md_pad_o_from_the_igor_mac),
      .md_padoe_o_from_the_igor_mac   (md_padoe_o_from_the_igor_mac),
      .mdc_pad_o_from_the_igor_mac    (mdc_pad_o_from_the_igor_mac),
      .mem_addr_from_the_ram          (mem_addr_from_the_ram),
      .mem_ba_from_the_ram            (mem_ba_from_the_ram),
      .mem_cas_n_from_the_ram         (mem_cas_n_from_the_ram),
      .mem_cke_from_the_ram           (mem_cke_from_the_ram),
      .mem_clk_n_to_and_from_the_ram  (mem_clk_n_to_and_from_the_ram),
      .mem_clk_to_and_from_the_ram    (mem_clk_to_and_from_the_ram),
      .mem_cs_n_from_the_ram          (mem_cs_n_from_the_ram),
      .mem_dm_from_the_ram            (mem_dm_from_the_ram),
      .mem_dq_to_and_from_the_ram     (mem_dq_to_and_from_the_ram),
      .mem_dqs_to_and_from_the_ram    (mem_dqs_to_and_from_the_ram),
      .mem_odt_from_the_ram           (mem_odt_from_the_ram),
      .mem_ras_n_from_the_ram         (mem_ras_n_from_the_ram),
      .mem_we_n_from_the_ram          (mem_we_n_from_the_ram),
      .mrx_clk_pad_i_to_the_igor_mac  (mrx_clk_pad_i_to_the_igor_mac),
      .mrxd_pad_i_to_the_igor_mac     (mrxd_pad_i_to_the_igor_mac),
      .mrxdv_pad_i_to_the_igor_mac    (mrxdv_pad_i_to_the_igor_mac),
      .mrxerr_pad_i_to_the_igor_mac   (mrxerr_pad_i_to_the_igor_mac),
      .mtx_clk_pad_i_to_the_igor_mac  (mtx_clk_pad_i_to_the_igor_mac),
      .mtxd_pad_o_from_the_igor_mac   (mtxd_pad_o_from_the_igor_mac),
      .mtxen_pad_o_from_the_igor_mac  (mtxen_pad_o_from_the_igor_mac),
      .mtxerr_pad_o_from_the_igor_mac (mtxerr_pad_o_from_the_igor_mac),
      .out_data_from_the_tx_table     (out_data_from_the_tx_table),
      .out_sync_from_the_tx_table     (out_sync_from_the_tx_table),
      .out_valid_from_the_tx_table    (out_valid_from_the_tx_table),
      .ram_aux_full_rate_clk_out      (ram_aux_full_rate_clk_out),
      .ram_aux_half_rate_clk_out      (ram_aux_half_rate_clk_out),
      .ram_phy_clk_out                (ram_phy_clk_out),
      .reset_n                        (reset_n),
      .reset_phy_clk_n_from_the_ram   (reset_phy_clk_n_from_the_ram),
      .rxd_to_the_uart_0              (rxd_to_the_uart_0),
      .sce_from_the_epcs_controller   (sce_from_the_epcs_controller),
      .sdo_from_the_epcs_controller   (sdo_from_the_epcs_controller),
      .txd_from_the_uart_0            (txd_from_the_uart_0)
    );

  initial
    clk_125 = 1'b0;
  always
    #4 clk_125 <= ~clk_125;
  
  initial 
    begin
      reset_n <= 0;
      #80 reset_n <= 1;
    end

endmodule


//synthesis translate_on