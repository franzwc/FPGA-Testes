


	

		
